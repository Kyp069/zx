//-------------------------------------------------------------------------------------------------
module mmcm1
//-------------------------------------------------------------------------------------------------
(
	input  wire ci,
	output wire co1,
	output wire locked
);
//-------------------------------------------------------------------------------------------------

wire fi1, fo1;

MMCME2_BASE #
(
	.CLKIN1_PERIOD   (20.000),
	.DIVCLK_DIVIDE   ( 3    ),
	.CLKFBOUT_MULT_F (51.500),
	.CLKOUT0_DIVIDE_F(15.125)
)
mmcm1
(
	.CLKIN1          (ci),
	.CLKFBIN         (fi1),

	.PWRDWN          (1'b0),
	.RST             (1'b0),

	.CLKFBOUT        (fo1),
	.CLKFBOUTB       (),
	.CLKOUT0         (co1),
	.CLKOUT0B        (),
	.CLKOUT1         (),
	.CLKOUT1B        (),
	.CLKOUT2         (),
	.CLKOUT2B        (),
	.CLKOUT3         (),
	.CLKOUT3B        (),
	.CLKOUT4         (),
	.CLKOUT5         (),
	.CLKOUT6         (),
	.LOCKED          (locked)
);

BUFG bufgfb1(.I(fo1), .O(fi1));

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
