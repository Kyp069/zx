//-------------------------------------------------------------------------------------------------
module flash
//-------------------------------------------------------------------------------------------------
(
	input  wire clock,

	output reg  vga,

	output reg  cs,
	output wire ck,
	output wire mosi,
	input  wire miso
);
//-------------------------------------------------------------------------------------------------

reg[3:0] ce = 0;
always @(negedge clock) ce <= ce+1'd1;

wire pe = ~ce[0] & ~ce[1] & ~ce[2] &  ce[3];
wire ne = ~ce[0] & ~ce[1] & ~ce[2];

//-------------------------------------------------------------------------------------------------

reg io;

reg[7:0] d;
reg[7:0] fc = 0;

always @(posedge clock) if(pe)
if(!fc[7]) begin
	fc <= fc+1'd1;

	case(fc)
		 0: cs <= 1'b1;
		14: cs <= 1'b0;

//		 0: begin tx <= 1'b1; d <= 8'h13; end
//		 1: begin tx <= 1'b0; end

		16: begin io <= 1'b1; d <= 8'h03; end // 8'h03
		17: begin io <= 1'b0; end

		32: begin io <= 1'b1; d <= 8'h00; end
		33: begin io <= 1'b0; end

		48: begin io <= 1'b1; d <= 8'h8F; end // 8'h70
		49: begin io <= 1'b0; end

		64: begin io <= 1'b1; d <= 8'hD5; end // 8'h4D
		65: begin io <= 1'b0; end

//		80: io <= 1'b1;
//		81: io <= 1'b0;

		96: begin io <= 1'b1; d <= 8'hFF; end
		97: begin io <= 1'b0; end

		98: vga <= q[1:0] == 2'b10;
		99: cs <= 1'b1;
	endcase
end

//-------------------------------------------------------------------------------------------------

wire[7:0] q;

spi Flash
(
	.clock  (clock  ),
	.ce     (ne     ),
	.io     (io     ),
	.d      (d      ),
	.q      (q      ),
	.ck     (ck     ),
	.mosi   (mosi   ),
	.miso   (miso   )
);

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
