
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c0",x"fb",x"c1",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c0",x"fb",x"c1"),
    14 => (x"48",x"ec",x"e9",x"c1"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c0",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e7",x"f8"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"72",x"1e",x"73"),
    21 => (x"ca",x"04",x"8b",x"c1"),
    22 => (x"11",x"48",x"12",x"87"),
    23 => (x"88",x"87",x"c4",x"02"),
    24 => (x"26",x"87",x"f1",x"02"),
    25 => (x"26",x"4b",x"26",x"4a"),
    26 => (x"48",x"73",x"1e",x"4f"),
    27 => (x"02",x"a9",x"73",x"81"),
    28 => (x"53",x"12",x"87",x"c5"),
    29 => (x"26",x"87",x"f6",x"05"),
    30 => (x"4a",x"71",x"1e",x"4f"),
    31 => (x"48",x"49",x"66",x"c4"),
    32 => (x"a6",x"c8",x"88",x"c1"),
    33 => (x"02",x"99",x"71",x"58"),
    34 => (x"d4",x"ff",x"87",x"d6"),
    35 => (x"78",x"ff",x"c3",x"48"),
    36 => (x"66",x"c4",x"52",x"68"),
    37 => (x"88",x"c1",x"48",x"49"),
    38 => (x"71",x"58",x"a6",x"c8"),
    39 => (x"87",x"ea",x"05",x"99"),
    40 => (x"73",x"1e",x"4f",x"26"),
    41 => (x"4b",x"d4",x"ff",x"1e"),
    42 => (x"6b",x"7b",x"ff",x"c3"),
    43 => (x"7b",x"ff",x"c3",x"4a"),
    44 => (x"32",x"c8",x"49",x"6b"),
    45 => (x"ff",x"c3",x"b1",x"72"),
    46 => (x"c8",x"4a",x"6b",x"7b"),
    47 => (x"c3",x"b2",x"71",x"31"),
    48 => (x"49",x"6b",x"7b",x"ff"),
    49 => (x"b1",x"72",x"32",x"c8"),
    50 => (x"87",x"c4",x"48",x"71"),
    51 => (x"4c",x"26",x"4d",x"26"),
    52 => (x"4f",x"26",x"4b",x"26"),
    53 => (x"5c",x"5b",x"5e",x"0e"),
    54 => (x"4a",x"71",x"0e",x"5d"),
    55 => (x"72",x"4c",x"d4",x"ff"),
    56 => (x"99",x"ff",x"c3",x"49"),
    57 => (x"e9",x"c1",x"7c",x"71"),
    58 => (x"c8",x"05",x"bf",x"ec"),
    59 => (x"48",x"66",x"d0",x"87"),
    60 => (x"a6",x"d4",x"30",x"c9"),
    61 => (x"49",x"66",x"d0",x"58"),
    62 => (x"ff",x"c3",x"29",x"d8"),
    63 => (x"d0",x"7c",x"71",x"99"),
    64 => (x"29",x"d0",x"49",x"66"),
    65 => (x"71",x"99",x"ff",x"c3"),
    66 => (x"49",x"66",x"d0",x"7c"),
    67 => (x"ff",x"c3",x"29",x"c8"),
    68 => (x"d0",x"7c",x"71",x"99"),
    69 => (x"ff",x"c3",x"49",x"66"),
    70 => (x"72",x"7c",x"71",x"99"),
    71 => (x"c3",x"29",x"d0",x"49"),
    72 => (x"7c",x"71",x"99",x"ff"),
    73 => (x"f0",x"c9",x"4b",x"6c"),
    74 => (x"ff",x"c3",x"4d",x"ff"),
    75 => (x"87",x"d0",x"05",x"ab"),
    76 => (x"6c",x"7c",x"ff",x"c3"),
    77 => (x"02",x"8d",x"c1",x"4b"),
    78 => (x"ff",x"c3",x"87",x"c6"),
    79 => (x"87",x"f0",x"02",x"ab"),
    80 => (x"c7",x"fe",x"48",x"73"),
    81 => (x"5b",x"5e",x"0e",x"87"),
    82 => (x"71",x"0e",x"5d",x"5c"),
    83 => (x"c5",x"4c",x"c0",x"4b"),
    84 => (x"4a",x"df",x"cd",x"ee"),
    85 => (x"c3",x"48",x"d4",x"ff"),
    86 => (x"49",x"68",x"78",x"ff"),
    87 => (x"05",x"a9",x"fe",x"c3"),
    88 => (x"70",x"87",x"fd",x"c0"),
    89 => (x"02",x"9b",x"73",x"4d"),
    90 => (x"66",x"d0",x"87",x"cc"),
    91 => (x"fc",x"49",x"73",x"1e"),
    92 => (x"86",x"c4",x"87",x"c7"),
    93 => (x"d0",x"ff",x"87",x"d6"),
    94 => (x"78",x"d1",x"c4",x"48"),
    95 => (x"d0",x"7d",x"ff",x"c3"),
    96 => (x"88",x"c1",x"48",x"66"),
    97 => (x"70",x"58",x"a6",x"d4"),
    98 => (x"87",x"f0",x"05",x"98"),
    99 => (x"c3",x"48",x"d4",x"ff"),
   100 => (x"73",x"78",x"78",x"ff"),
   101 => (x"87",x"c5",x"05",x"9b"),
   102 => (x"d0",x"48",x"d0",x"ff"),
   103 => (x"4c",x"4a",x"c1",x"78"),
   104 => (x"fe",x"05",x"8a",x"c1"),
   105 => (x"48",x"74",x"87",x"ee"),
   106 => (x"1e",x"87",x"e1",x"fc"),
   107 => (x"4a",x"71",x"1e",x"73"),
   108 => (x"d4",x"ff",x"4b",x"c0"),
   109 => (x"78",x"ff",x"c3",x"48"),
   110 => (x"c4",x"48",x"d0",x"ff"),
   111 => (x"d4",x"ff",x"78",x"c3"),
   112 => (x"78",x"ff",x"c3",x"48"),
   113 => (x"ff",x"c0",x"1e",x"72"),
   114 => (x"49",x"d1",x"c1",x"f0"),
   115 => (x"c4",x"87",x"c5",x"fc"),
   116 => (x"05",x"98",x"70",x"86"),
   117 => (x"c0",x"c8",x"87",x"d2"),
   118 => (x"49",x"66",x"cc",x"1e"),
   119 => (x"c4",x"87",x"e6",x"fd"),
   120 => (x"ff",x"4b",x"70",x"86"),
   121 => (x"78",x"c2",x"48",x"d0"),
   122 => (x"e3",x"fb",x"48",x"73"),
   123 => (x"5b",x"5e",x"0e",x"87"),
   124 => (x"f8",x"0e",x"5d",x"5c"),
   125 => (x"c4",x"f2",x"c1",x"86"),
   126 => (x"c1",x"78",x"c0",x"48"),
   127 => (x"c0",x"1e",x"fc",x"e9"),
   128 => (x"87",x"e7",x"fe",x"49"),
   129 => (x"98",x"70",x"86",x"c4"),
   130 => (x"c0",x"87",x"c5",x"05"),
   131 => (x"87",x"c7",x"c9",x"48"),
   132 => (x"7e",x"c1",x"4d",x"c0"),
   133 => (x"49",x"bf",x"ec",x"da"),
   134 => (x"4a",x"f2",x"ea",x"c1"),
   135 => (x"f8",x"4b",x"c8",x"71"),
   136 => (x"98",x"70",x"87",x"ed"),
   137 => (x"c0",x"87",x"c2",x"05"),
   138 => (x"bf",x"e8",x"da",x"7e"),
   139 => (x"ce",x"eb",x"c1",x"49"),
   140 => (x"4b",x"c8",x"71",x"4a"),
   141 => (x"70",x"87",x"d8",x"f8"),
   142 => (x"87",x"c2",x"05",x"98"),
   143 => (x"02",x"6e",x"7e",x"c0"),
   144 => (x"c1",x"87",x"fd",x"c0"),
   145 => (x"4d",x"bf",x"c2",x"f1"),
   146 => (x"9f",x"fa",x"f1",x"c1"),
   147 => (x"c5",x"48",x"7e",x"bf"),
   148 => (x"05",x"a8",x"ea",x"d6"),
   149 => (x"f1",x"c1",x"87",x"c7"),
   150 => (x"ce",x"4d",x"bf",x"c2"),
   151 => (x"ca",x"48",x"6e",x"87"),
   152 => (x"02",x"a8",x"d5",x"e9"),
   153 => (x"48",x"c0",x"87",x"c5"),
   154 => (x"c1",x"87",x"ec",x"c7"),
   155 => (x"75",x"1e",x"fc",x"e9"),
   156 => (x"87",x"f7",x"fc",x"49"),
   157 => (x"98",x"70",x"86",x"c4"),
   158 => (x"c0",x"87",x"c5",x"05"),
   159 => (x"87",x"d7",x"c7",x"48"),
   160 => (x"49",x"bf",x"e8",x"da"),
   161 => (x"4a",x"ce",x"eb",x"c1"),
   162 => (x"f7",x"4b",x"c8",x"71"),
   163 => (x"98",x"70",x"87",x"c1"),
   164 => (x"c1",x"87",x"c8",x"05"),
   165 => (x"c1",x"48",x"c4",x"f2"),
   166 => (x"da",x"87",x"d8",x"78"),
   167 => (x"c1",x"49",x"bf",x"ec"),
   168 => (x"71",x"4a",x"f2",x"ea"),
   169 => (x"e6",x"f6",x"4b",x"c8"),
   170 => (x"02",x"98",x"70",x"87"),
   171 => (x"48",x"c0",x"87",x"c5"),
   172 => (x"c1",x"87",x"e4",x"c6"),
   173 => (x"bf",x"97",x"fa",x"f1"),
   174 => (x"a9",x"d5",x"c1",x"49"),
   175 => (x"c1",x"87",x"cd",x"05"),
   176 => (x"bf",x"97",x"fb",x"f1"),
   177 => (x"a9",x"ea",x"c2",x"49"),
   178 => (x"87",x"c5",x"c0",x"02"),
   179 => (x"c6",x"c6",x"48",x"c0"),
   180 => (x"fc",x"e9",x"c1",x"87"),
   181 => (x"48",x"7e",x"bf",x"97"),
   182 => (x"02",x"a8",x"e9",x"c3"),
   183 => (x"6e",x"87",x"ce",x"c0"),
   184 => (x"a8",x"eb",x"c3",x"48"),
   185 => (x"87",x"c5",x"c0",x"02"),
   186 => (x"ea",x"c5",x"48",x"c0"),
   187 => (x"c7",x"ea",x"c1",x"87"),
   188 => (x"99",x"49",x"bf",x"97"),
   189 => (x"87",x"cc",x"c0",x"05"),
   190 => (x"97",x"c8",x"ea",x"c1"),
   191 => (x"a9",x"c2",x"49",x"bf"),
   192 => (x"87",x"c5",x"c0",x"02"),
   193 => (x"ce",x"c5",x"48",x"c0"),
   194 => (x"c9",x"ea",x"c1",x"87"),
   195 => (x"c1",x"48",x"bf",x"97"),
   196 => (x"70",x"58",x"c0",x"f2"),
   197 => (x"88",x"c1",x"48",x"4c"),
   198 => (x"58",x"c4",x"f2",x"c1"),
   199 => (x"97",x"ca",x"ea",x"c1"),
   200 => (x"81",x"75",x"49",x"bf"),
   201 => (x"97",x"cb",x"ea",x"c1"),
   202 => (x"32",x"c8",x"4a",x"bf"),
   203 => (x"c1",x"7e",x"a1",x"72"),
   204 => (x"6e",x"48",x"d1",x"f6"),
   205 => (x"cc",x"ea",x"c1",x"78"),
   206 => (x"c8",x"48",x"bf",x"97"),
   207 => (x"f2",x"c1",x"58",x"a6"),
   208 => (x"c2",x"02",x"bf",x"c4"),
   209 => (x"e8",x"da",x"87",x"d3"),
   210 => (x"eb",x"c1",x"49",x"bf"),
   211 => (x"c8",x"71",x"4a",x"ce"),
   212 => (x"87",x"fb",x"f3",x"4b"),
   213 => (x"c0",x"02",x"98",x"70"),
   214 => (x"48",x"c0",x"87",x"c5"),
   215 => (x"c1",x"87",x"f8",x"c3"),
   216 => (x"4c",x"bf",x"fc",x"f1"),
   217 => (x"5c",x"e5",x"f6",x"c1"),
   218 => (x"97",x"e1",x"ea",x"c1"),
   219 => (x"31",x"c8",x"49",x"bf"),
   220 => (x"97",x"e0",x"ea",x"c1"),
   221 => (x"49",x"a1",x"4a",x"bf"),
   222 => (x"97",x"e2",x"ea",x"c1"),
   223 => (x"32",x"d0",x"4a",x"bf"),
   224 => (x"c1",x"49",x"a1",x"72"),
   225 => (x"bf",x"97",x"e3",x"ea"),
   226 => (x"72",x"32",x"d8",x"4a"),
   227 => (x"66",x"c4",x"49",x"a1"),
   228 => (x"d1",x"f6",x"c1",x"91"),
   229 => (x"f6",x"c1",x"81",x"bf"),
   230 => (x"ea",x"c1",x"59",x"d9"),
   231 => (x"4a",x"bf",x"97",x"e9"),
   232 => (x"ea",x"c1",x"32",x"c8"),
   233 => (x"4b",x"bf",x"97",x"e8"),
   234 => (x"ea",x"c1",x"4a",x"a2"),
   235 => (x"4b",x"bf",x"97",x"ea"),
   236 => (x"a2",x"73",x"33",x"d0"),
   237 => (x"eb",x"ea",x"c1",x"4a"),
   238 => (x"cf",x"4b",x"bf",x"97"),
   239 => (x"73",x"33",x"d8",x"9b"),
   240 => (x"f6",x"c1",x"4a",x"a2"),
   241 => (x"f6",x"c1",x"5a",x"dd"),
   242 => (x"c2",x"4a",x"bf",x"d9"),
   243 => (x"c1",x"92",x"74",x"8a"),
   244 => (x"72",x"48",x"dd",x"f6"),
   245 => (x"ca",x"c1",x"78",x"a1"),
   246 => (x"ce",x"ea",x"c1",x"87"),
   247 => (x"c8",x"49",x"bf",x"97"),
   248 => (x"cd",x"ea",x"c1",x"31"),
   249 => (x"a1",x"4a",x"bf",x"97"),
   250 => (x"cc",x"f2",x"c1",x"49"),
   251 => (x"c8",x"f2",x"c1",x"59"),
   252 => (x"31",x"c5",x"49",x"bf"),
   253 => (x"c9",x"81",x"ff",x"c7"),
   254 => (x"e5",x"f6",x"c1",x"29"),
   255 => (x"d3",x"ea",x"c1",x"59"),
   256 => (x"c8",x"4a",x"bf",x"97"),
   257 => (x"d2",x"ea",x"c1",x"32"),
   258 => (x"a2",x"4b",x"bf",x"97"),
   259 => (x"92",x"66",x"c4",x"4a"),
   260 => (x"f6",x"c1",x"82",x"6e"),
   261 => (x"f6",x"c1",x"5a",x"e1"),
   262 => (x"78",x"c0",x"48",x"d9"),
   263 => (x"48",x"d5",x"f6",x"c1"),
   264 => (x"c1",x"78",x"a1",x"72"),
   265 => (x"c1",x"48",x"e5",x"f6"),
   266 => (x"78",x"bf",x"d9",x"f6"),
   267 => (x"48",x"e9",x"f6",x"c1"),
   268 => (x"bf",x"dd",x"f6",x"c1"),
   269 => (x"c4",x"f2",x"c1",x"78"),
   270 => (x"c9",x"c0",x"02",x"bf"),
   271 => (x"c4",x"48",x"74",x"87"),
   272 => (x"c0",x"7e",x"70",x"30"),
   273 => (x"f6",x"c1",x"87",x"c9"),
   274 => (x"c4",x"48",x"bf",x"e1"),
   275 => (x"c1",x"7e",x"70",x"30"),
   276 => (x"6e",x"48",x"c8",x"f2"),
   277 => (x"f8",x"48",x"c1",x"78"),
   278 => (x"26",x"4d",x"26",x"8e"),
   279 => (x"26",x"4b",x"26",x"4c"),
   280 => (x"5b",x"5e",x"0e",x"4f"),
   281 => (x"71",x"0e",x"5d",x"5c"),
   282 => (x"c4",x"f2",x"c1",x"4a"),
   283 => (x"87",x"cb",x"02",x"bf"),
   284 => (x"2b",x"c7",x"4b",x"72"),
   285 => (x"ff",x"c1",x"4c",x"72"),
   286 => (x"72",x"87",x"c9",x"9c"),
   287 => (x"72",x"2b",x"c8",x"4b"),
   288 => (x"9c",x"ff",x"c3",x"4c"),
   289 => (x"bf",x"d1",x"f6",x"c1"),
   290 => (x"bf",x"e4",x"da",x"83"),
   291 => (x"87",x"d8",x"02",x"ab"),
   292 => (x"c1",x"5b",x"e8",x"da"),
   293 => (x"73",x"1e",x"fc",x"e9"),
   294 => (x"87",x"cf",x"f4",x"49"),
   295 => (x"98",x"70",x"86",x"c4"),
   296 => (x"c0",x"87",x"c5",x"05"),
   297 => (x"87",x"e6",x"c0",x"48"),
   298 => (x"bf",x"c4",x"f2",x"c1"),
   299 => (x"74",x"87",x"d2",x"02"),
   300 => (x"c1",x"91",x"c4",x"49"),
   301 => (x"69",x"81",x"fc",x"e9"),
   302 => (x"ff",x"ff",x"cf",x"4d"),
   303 => (x"cb",x"9d",x"ff",x"ff"),
   304 => (x"c2",x"49",x"74",x"87"),
   305 => (x"fc",x"e9",x"c1",x"91"),
   306 => (x"4d",x"69",x"9f",x"81"),
   307 => (x"c8",x"fe",x"48",x"75"),
   308 => (x"5b",x"5e",x"0e",x"87"),
   309 => (x"f4",x"0e",x"5d",x"5c"),
   310 => (x"c0",x"4a",x"71",x"86"),
   311 => (x"02",x"9a",x"72",x"7e"),
   312 => (x"e9",x"c1",x"87",x"d8"),
   313 => (x"78",x"c0",x"48",x"f8"),
   314 => (x"48",x"f0",x"e9",x"c1"),
   315 => (x"bf",x"e9",x"f6",x"c1"),
   316 => (x"f4",x"e9",x"c1",x"78"),
   317 => (x"e5",x"f6",x"c1",x"48"),
   318 => (x"f2",x"c1",x"78",x"bf"),
   319 => (x"50",x"c0",x"48",x"d9"),
   320 => (x"bf",x"c8",x"f2",x"c1"),
   321 => (x"f8",x"e9",x"c1",x"49"),
   322 => (x"aa",x"71",x"4a",x"bf"),
   323 => (x"87",x"c1",x"c4",x"03"),
   324 => (x"99",x"cf",x"49",x"72"),
   325 => (x"87",x"e7",x"c0",x"05"),
   326 => (x"c1",x"48",x"e4",x"da"),
   327 => (x"78",x"bf",x"f0",x"e9"),
   328 => (x"1e",x"fc",x"e9",x"c1"),
   329 => (x"bf",x"f0",x"e9",x"c1"),
   330 => (x"f0",x"e9",x"c1",x"49"),
   331 => (x"78",x"a1",x"c1",x"48"),
   332 => (x"87",x"f7",x"f1",x"71"),
   333 => (x"e0",x"da",x"86",x"c4"),
   334 => (x"fc",x"e9",x"c1",x"48"),
   335 => (x"da",x"87",x"ca",x"78"),
   336 => (x"c0",x"48",x"bf",x"e0"),
   337 => (x"e4",x"da",x"80",x"e0"),
   338 => (x"f8",x"e9",x"c1",x"58"),
   339 => (x"80",x"c1",x"48",x"bf"),
   340 => (x"58",x"fc",x"e9",x"c1"),
   341 => (x"00",x"06",x"a0",x"27"),
   342 => (x"bf",x"97",x"bf",x"00"),
   343 => (x"c2",x"02",x"9d",x"4d"),
   344 => (x"e5",x"c3",x"87",x"df"),
   345 => (x"d8",x"c2",x"02",x"ad"),
   346 => (x"bf",x"e0",x"da",x"87"),
   347 => (x"49",x"a3",x"cb",x"4b"),
   348 => (x"ac",x"cf",x"4c",x"11"),
   349 => (x"87",x"d2",x"c1",x"05"),
   350 => (x"99",x"df",x"49",x"75"),
   351 => (x"91",x"cd",x"89",x"c1"),
   352 => (x"81",x"cc",x"f2",x"c1"),
   353 => (x"12",x"4a",x"a3",x"c1"),
   354 => (x"4a",x"a3",x"c3",x"51"),
   355 => (x"a3",x"c5",x"51",x"12"),
   356 => (x"c7",x"51",x"12",x"4a"),
   357 => (x"51",x"12",x"4a",x"a3"),
   358 => (x"12",x"4a",x"a3",x"c9"),
   359 => (x"4a",x"a3",x"ce",x"51"),
   360 => (x"a3",x"d0",x"51",x"12"),
   361 => (x"d2",x"51",x"12",x"4a"),
   362 => (x"51",x"12",x"4a",x"a3"),
   363 => (x"12",x"4a",x"a3",x"d4"),
   364 => (x"4a",x"a3",x"d6",x"51"),
   365 => (x"a3",x"d8",x"51",x"12"),
   366 => (x"dc",x"51",x"12",x"4a"),
   367 => (x"51",x"12",x"4a",x"a3"),
   368 => (x"12",x"4a",x"a3",x"de"),
   369 => (x"c0",x"7e",x"c1",x"51"),
   370 => (x"49",x"74",x"87",x"f7"),
   371 => (x"c0",x"05",x"99",x"c8"),
   372 => (x"49",x"74",x"87",x"e8"),
   373 => (x"cf",x"05",x"99",x"d0"),
   374 => (x"02",x"66",x"dc",x"87"),
   375 => (x"49",x"73",x"87",x"ca"),
   376 => (x"70",x"0f",x"66",x"dc"),
   377 => (x"87",x"d2",x"02",x"98"),
   378 => (x"c6",x"c0",x"05",x"6e"),
   379 => (x"cc",x"f2",x"c1",x"87"),
   380 => (x"da",x"50",x"c0",x"48"),
   381 => (x"c2",x"48",x"bf",x"e0"),
   382 => (x"f2",x"c1",x"87",x"e1"),
   383 => (x"50",x"c0",x"48",x"d9"),
   384 => (x"c8",x"f2",x"c1",x"7e"),
   385 => (x"e9",x"c1",x"49",x"bf"),
   386 => (x"71",x"4a",x"bf",x"f8"),
   387 => (x"ff",x"fb",x"04",x"aa"),
   388 => (x"e9",x"f6",x"c1",x"87"),
   389 => (x"c8",x"c0",x"05",x"bf"),
   390 => (x"c4",x"f2",x"c1",x"87"),
   391 => (x"f8",x"c1",x"02",x"bf"),
   392 => (x"f4",x"e9",x"c1",x"87"),
   393 => (x"f8",x"f8",x"49",x"bf"),
   394 => (x"c1",x"49",x"70",x"87"),
   395 => (x"c4",x"59",x"f8",x"e9"),
   396 => (x"e9",x"c1",x"48",x"a6"),
   397 => (x"c1",x"78",x"bf",x"f4"),
   398 => (x"02",x"bf",x"c4",x"f2"),
   399 => (x"c4",x"87",x"d8",x"c0"),
   400 => (x"ff",x"cf",x"49",x"66"),
   401 => (x"99",x"f8",x"ff",x"ff"),
   402 => (x"c5",x"c0",x"02",x"a9"),
   403 => (x"c0",x"4c",x"c0",x"87"),
   404 => (x"4c",x"c1",x"87",x"e1"),
   405 => (x"c4",x"87",x"dc",x"c0"),
   406 => (x"ff",x"cf",x"49",x"66"),
   407 => (x"02",x"a9",x"99",x"f8"),
   408 => (x"c8",x"87",x"c8",x"c0"),
   409 => (x"78",x"c0",x"48",x"a6"),
   410 => (x"c8",x"87",x"c5",x"c0"),
   411 => (x"78",x"c1",x"48",x"a6"),
   412 => (x"74",x"4c",x"66",x"c8"),
   413 => (x"e0",x"c0",x"05",x"9c"),
   414 => (x"49",x"66",x"c4",x"87"),
   415 => (x"f1",x"c1",x"89",x"c2"),
   416 => (x"91",x"4a",x"bf",x"fc"),
   417 => (x"bf",x"d5",x"f6",x"c1"),
   418 => (x"f0",x"e9",x"c1",x"4a"),
   419 => (x"78",x"a1",x"72",x"48"),
   420 => (x"48",x"f8",x"e9",x"c1"),
   421 => (x"e7",x"f9",x"78",x"c0"),
   422 => (x"f4",x"48",x"c0",x"87"),
   423 => (x"87",x"f9",x"f6",x"8e"),
   424 => (x"00",x"00",x"00",x"00"),
   425 => (x"ff",x"ff",x"ff",x"ff"),
   426 => (x"00",x"00",x"06",x"b0"),
   427 => (x"00",x"00",x"06",x"b9"),
   428 => (x"33",x"54",x"41",x"46"),
   429 => (x"20",x"20",x"20",x"32"),
   430 => (x"54",x"41",x"46",x"00"),
   431 => (x"20",x"20",x"36",x"31"),
   432 => (x"ff",x"1e",x"00",x"20"),
   433 => (x"ff",x"c3",x"48",x"d4"),
   434 => (x"26",x"48",x"68",x"78"),
   435 => (x"d4",x"ff",x"1e",x"4f"),
   436 => (x"78",x"ff",x"c3",x"48"),
   437 => (x"c0",x"48",x"d0",x"ff"),
   438 => (x"d4",x"ff",x"78",x"e1"),
   439 => (x"c1",x"78",x"d4",x"48"),
   440 => (x"ff",x"48",x"ed",x"f6"),
   441 => (x"26",x"50",x"bf",x"d4"),
   442 => (x"d0",x"ff",x"1e",x"4f"),
   443 => (x"78",x"e0",x"c0",x"48"),
   444 => (x"ff",x"1e",x"4f",x"26"),
   445 => (x"49",x"70",x"87",x"cc"),
   446 => (x"87",x"c6",x"02",x"99"),
   447 => (x"05",x"a9",x"fb",x"c0"),
   448 => (x"48",x"71",x"87",x"f1"),
   449 => (x"5e",x"0e",x"4f",x"26"),
   450 => (x"71",x"0e",x"5c",x"5b"),
   451 => (x"fe",x"4c",x"c0",x"4b"),
   452 => (x"49",x"70",x"87",x"f0"),
   453 => (x"f9",x"c0",x"02",x"99"),
   454 => (x"a9",x"ec",x"c0",x"87"),
   455 => (x"87",x"f2",x"c0",x"02"),
   456 => (x"02",x"a9",x"fb",x"c0"),
   457 => (x"cc",x"87",x"eb",x"c0"),
   458 => (x"03",x"ac",x"b7",x"66"),
   459 => (x"66",x"d0",x"87",x"c7"),
   460 => (x"71",x"87",x"c2",x"02"),
   461 => (x"02",x"99",x"71",x"53"),
   462 => (x"84",x"c1",x"87",x"c2"),
   463 => (x"70",x"87",x"c3",x"fe"),
   464 => (x"cd",x"02",x"99",x"49"),
   465 => (x"a9",x"ec",x"c0",x"87"),
   466 => (x"c0",x"87",x"c7",x"02"),
   467 => (x"ff",x"05",x"a9",x"fb"),
   468 => (x"66",x"d0",x"87",x"d5"),
   469 => (x"c0",x"87",x"c3",x"02"),
   470 => (x"ec",x"c0",x"7b",x"97"),
   471 => (x"87",x"c4",x"05",x"a9"),
   472 => (x"87",x"c5",x"4a",x"74"),
   473 => (x"0a",x"c0",x"4a",x"74"),
   474 => (x"c2",x"48",x"72",x"8a"),
   475 => (x"26",x"4d",x"26",x"87"),
   476 => (x"26",x"4b",x"26",x"4c"),
   477 => (x"c9",x"fd",x"1e",x"4f"),
   478 => (x"4a",x"49",x"70",x"87"),
   479 => (x"04",x"aa",x"f0",x"c0"),
   480 => (x"f9",x"c0",x"87",x"c9"),
   481 => (x"87",x"c3",x"01",x"aa"),
   482 => (x"c1",x"8a",x"f0",x"c0"),
   483 => (x"c9",x"04",x"aa",x"c1"),
   484 => (x"aa",x"da",x"c1",x"87"),
   485 => (x"c0",x"87",x"c3",x"01"),
   486 => (x"48",x"72",x"8a",x"f7"),
   487 => (x"5e",x"0e",x"4f",x"26"),
   488 => (x"0e",x"5d",x"5c",x"5b"),
   489 => (x"4c",x"71",x"86",x"f8"),
   490 => (x"e0",x"fc",x"7e",x"c0"),
   491 => (x"c0",x"4b",x"c0",x"87"),
   492 => (x"bf",x"97",x"cb",x"e1"),
   493 => (x"04",x"a9",x"c0",x"49"),
   494 => (x"f5",x"fc",x"87",x"cf"),
   495 => (x"c0",x"83",x"c1",x"87"),
   496 => (x"bf",x"97",x"cb",x"e1"),
   497 => (x"f1",x"06",x"ab",x"49"),
   498 => (x"cb",x"e1",x"c0",x"87"),
   499 => (x"cf",x"02",x"bf",x"97"),
   500 => (x"87",x"ee",x"fb",x"87"),
   501 => (x"02",x"99",x"49",x"70"),
   502 => (x"ec",x"c0",x"87",x"c6"),
   503 => (x"87",x"f1",x"05",x"a9"),
   504 => (x"dd",x"fb",x"4b",x"c0"),
   505 => (x"fb",x"4d",x"70",x"87"),
   506 => (x"a6",x"c8",x"87",x"d8"),
   507 => (x"87",x"d2",x"fb",x"58"),
   508 => (x"83",x"c1",x"4a",x"70"),
   509 => (x"97",x"49",x"a4",x"c8"),
   510 => (x"02",x"ad",x"49",x"69"),
   511 => (x"ff",x"c0",x"87",x"c7"),
   512 => (x"e7",x"c0",x"05",x"ad"),
   513 => (x"49",x"a4",x"c9",x"87"),
   514 => (x"c4",x"49",x"69",x"97"),
   515 => (x"c7",x"02",x"a9",x"66"),
   516 => (x"ff",x"c0",x"48",x"87"),
   517 => (x"87",x"d4",x"05",x"a8"),
   518 => (x"97",x"49",x"a4",x"ca"),
   519 => (x"02",x"aa",x"49",x"69"),
   520 => (x"ff",x"c0",x"87",x"c6"),
   521 => (x"87",x"c4",x"05",x"aa"),
   522 => (x"87",x"d0",x"7e",x"c1"),
   523 => (x"02",x"ad",x"ec",x"c0"),
   524 => (x"fb",x"c0",x"87",x"c6"),
   525 => (x"87",x"c4",x"05",x"ad"),
   526 => (x"7e",x"c1",x"4b",x"c0"),
   527 => (x"e1",x"fe",x"02",x"6e"),
   528 => (x"87",x"e5",x"fa",x"87"),
   529 => (x"8e",x"f8",x"48",x"73"),
   530 => (x"00",x"87",x"e2",x"fc"),
   531 => (x"5c",x"5b",x"5e",x"0e"),
   532 => (x"71",x"1e",x"0e",x"5d"),
   533 => (x"4d",x"4c",x"c0",x"4b"),
   534 => (x"e7",x"c0",x"04",x"ab"),
   535 => (x"1e",x"de",x"de",x"87"),
   536 => (x"c4",x"02",x"9d",x"75"),
   537 => (x"c2",x"4a",x"c0",x"87"),
   538 => (x"72",x"4a",x"c1",x"87"),
   539 => (x"87",x"e1",x"f1",x"49"),
   540 => (x"7e",x"70",x"86",x"c4"),
   541 => (x"05",x"6e",x"84",x"c1"),
   542 => (x"4c",x"73",x"87",x"c2"),
   543 => (x"ac",x"73",x"85",x"c1"),
   544 => (x"87",x"d9",x"ff",x"06"),
   545 => (x"26",x"26",x"48",x"6e"),
   546 => (x"26",x"4c",x"26",x"4d"),
   547 => (x"1e",x"4f",x"26",x"4b"),
   548 => (x"c0",x"1e",x"4f",x"26"),
   549 => (x"1e",x"4f",x"26",x"48"),
   550 => (x"cb",x"49",x"4a",x"71"),
   551 => (x"d6",x"fa",x"c0",x"91"),
   552 => (x"11",x"81",x"c8",x"81"),
   553 => (x"f2",x"f6",x"c1",x"48"),
   554 => (x"f2",x"f6",x"c1",x"58"),
   555 => (x"c1",x"78",x"c0",x"48"),
   556 => (x"87",x"ea",x"d5",x"49"),
   557 => (x"c0",x"1e",x"4f",x"26"),
   558 => (x"d2",x"f9",x"c0",x"49"),
   559 => (x"1e",x"4f",x"26",x"87"),
   560 => (x"d2",x"02",x"99",x"71"),
   561 => (x"eb",x"fb",x"c0",x"87"),
   562 => (x"f7",x"50",x"c0",x"48"),
   563 => (x"d7",x"e2",x"c0",x"80"),
   564 => (x"cf",x"fa",x"c0",x"40"),
   565 => (x"c0",x"87",x"ce",x"78"),
   566 => (x"c0",x"48",x"e7",x"fb"),
   567 => (x"fc",x"78",x"c8",x"fa"),
   568 => (x"f6",x"e2",x"c0",x"80"),
   569 => (x"0e",x"4f",x"26",x"78"),
   570 => (x"0e",x"5c",x"5b",x"5e"),
   571 => (x"cb",x"4a",x"4c",x"71"),
   572 => (x"d6",x"fa",x"c0",x"92"),
   573 => (x"49",x"a2",x"c8",x"82"),
   574 => (x"97",x"4b",x"a2",x"c9"),
   575 => (x"97",x"1e",x"4b",x"6b"),
   576 => (x"ca",x"1e",x"49",x"69"),
   577 => (x"c0",x"49",x"12",x"82"),
   578 => (x"c0",x"87",x"cd",x"e4"),
   579 => (x"87",x"ce",x"d4",x"49"),
   580 => (x"f6",x"c0",x"49",x"74"),
   581 => (x"8e",x"f8",x"87",x"d4"),
   582 => (x"1e",x"87",x"ee",x"fd"),
   583 => (x"4b",x"71",x"1e",x"73"),
   584 => (x"87",x"c3",x"ff",x"49"),
   585 => (x"fe",x"fe",x"49",x"73"),
   586 => (x"c0",x"49",x"c0",x"87"),
   587 => (x"fd",x"87",x"e0",x"f7"),
   588 => (x"73",x"1e",x"87",x"d9"),
   589 => (x"c6",x"4b",x"71",x"1e"),
   590 => (x"db",x"02",x"4a",x"a3"),
   591 => (x"02",x"8a",x"c1",x"87"),
   592 => (x"02",x"8a",x"87",x"d6"),
   593 => (x"8a",x"87",x"da",x"c1"),
   594 => (x"87",x"fc",x"c0",x"02"),
   595 => (x"e1",x"c0",x"02",x"8a"),
   596 => (x"cb",x"02",x"8a",x"87"),
   597 => (x"87",x"db",x"c1",x"87"),
   598 => (x"fa",x"fc",x"49",x"c7"),
   599 => (x"87",x"de",x"c1",x"87"),
   600 => (x"bf",x"f2",x"f6",x"c1"),
   601 => (x"87",x"cb",x"c1",x"02"),
   602 => (x"c1",x"88",x"c1",x"48"),
   603 => (x"c1",x"58",x"f6",x"f6"),
   604 => (x"f6",x"c1",x"87",x"c1"),
   605 => (x"c0",x"02",x"bf",x"f6"),
   606 => (x"f6",x"c1",x"87",x"f9"),
   607 => (x"c1",x"48",x"bf",x"f2"),
   608 => (x"f6",x"f6",x"c1",x"80"),
   609 => (x"87",x"eb",x"c0",x"58"),
   610 => (x"bf",x"f2",x"f6",x"c1"),
   611 => (x"c1",x"89",x"c6",x"49"),
   612 => (x"c0",x"59",x"f6",x"f6"),
   613 => (x"da",x"03",x"a9",x"b7"),
   614 => (x"f2",x"f6",x"c1",x"87"),
   615 => (x"d2",x"78",x"c0",x"48"),
   616 => (x"f6",x"f6",x"c1",x"87"),
   617 => (x"87",x"cb",x"02",x"bf"),
   618 => (x"bf",x"f2",x"f6",x"c1"),
   619 => (x"c1",x"80",x"c6",x"48"),
   620 => (x"c0",x"58",x"f6",x"f6"),
   621 => (x"87",x"e6",x"d1",x"49"),
   622 => (x"f3",x"c0",x"49",x"73"),
   623 => (x"ca",x"fb",x"87",x"ec"),
   624 => (x"5b",x"5e",x"0e",x"87"),
   625 => (x"ff",x"0e",x"5d",x"5c"),
   626 => (x"a6",x"dc",x"86",x"d0"),
   627 => (x"48",x"a6",x"c8",x"59"),
   628 => (x"80",x"c4",x"78",x"c0"),
   629 => (x"78",x"66",x"c4",x"c1"),
   630 => (x"78",x"c1",x"80",x"c4"),
   631 => (x"78",x"c1",x"80",x"c4"),
   632 => (x"48",x"f6",x"f6",x"c1"),
   633 => (x"f6",x"c1",x"78",x"c1"),
   634 => (x"de",x"48",x"bf",x"ee"),
   635 => (x"87",x"cb",x"05",x"a8"),
   636 => (x"70",x"87",x"df",x"fa"),
   637 => (x"59",x"a6",x"cc",x"49"),
   638 => (x"f3",x"87",x"e3",x"cf"),
   639 => (x"f1",x"f3",x"87",x"cf"),
   640 => (x"87",x"fe",x"f2",x"87"),
   641 => (x"fb",x"c0",x"4c",x"70"),
   642 => (x"fb",x"c1",x"02",x"ac"),
   643 => (x"05",x"66",x"d8",x"87"),
   644 => (x"c1",x"87",x"ed",x"c1"),
   645 => (x"c4",x"4a",x"66",x"c0"),
   646 => (x"72",x"7e",x"6a",x"82"),
   647 => (x"d2",x"f8",x"c0",x"1e"),
   648 => (x"49",x"66",x"c4",x"48"),
   649 => (x"20",x"4a",x"a1",x"c8"),
   650 => (x"05",x"aa",x"71",x"41"),
   651 => (x"51",x"10",x"87",x"f9"),
   652 => (x"c0",x"c1",x"4a",x"26"),
   653 => (x"e2",x"c0",x"48",x"66"),
   654 => (x"49",x"6a",x"78",x"cf"),
   655 => (x"51",x"74",x"81",x"c7"),
   656 => (x"49",x"66",x"c0",x"c1"),
   657 => (x"51",x"c1",x"81",x"c8"),
   658 => (x"49",x"66",x"c0",x"c1"),
   659 => (x"51",x"c0",x"81",x"c9"),
   660 => (x"49",x"66",x"c0",x"c1"),
   661 => (x"51",x"c0",x"81",x"ca"),
   662 => (x"1e",x"d8",x"1e",x"c1"),
   663 => (x"81",x"c8",x"49",x"6a"),
   664 => (x"c8",x"87",x"e3",x"f2"),
   665 => (x"66",x"c4",x"c1",x"86"),
   666 => (x"01",x"a8",x"c0",x"48"),
   667 => (x"a6",x"c8",x"87",x"c7"),
   668 => (x"ce",x"78",x"c1",x"48"),
   669 => (x"66",x"c4",x"c1",x"87"),
   670 => (x"d0",x"88",x"c1",x"48"),
   671 => (x"87",x"c3",x"58",x"a6"),
   672 => (x"d0",x"87",x"ef",x"f1"),
   673 => (x"78",x"c2",x"48",x"a6"),
   674 => (x"cd",x"02",x"9c",x"74"),
   675 => (x"66",x"c8",x"87",x"cd"),
   676 => (x"66",x"c8",x"c1",x"48"),
   677 => (x"c2",x"cd",x"03",x"a8"),
   678 => (x"48",x"a6",x"dc",x"87"),
   679 => (x"80",x"e8",x"78",x"c0"),
   680 => (x"dd",x"f0",x"78",x"c0"),
   681 => (x"c1",x"4c",x"70",x"87"),
   682 => (x"c2",x"05",x"ac",x"d0"),
   683 => (x"66",x"c4",x"87",x"d6"),
   684 => (x"87",x"c1",x"f3",x"7e"),
   685 => (x"a6",x"c8",x"49",x"70"),
   686 => (x"87",x"c6",x"f0",x"59"),
   687 => (x"ec",x"c0",x"4c",x"70"),
   688 => (x"ea",x"c1",x"05",x"ac"),
   689 => (x"49",x"66",x"c8",x"87"),
   690 => (x"c0",x"c1",x"91",x"cb"),
   691 => (x"a1",x"c4",x"81",x"66"),
   692 => (x"c8",x"4d",x"6a",x"4a"),
   693 => (x"66",x"c4",x"4a",x"a1"),
   694 => (x"d7",x"e2",x"c0",x"52"),
   695 => (x"87",x"e2",x"ef",x"79"),
   696 => (x"02",x"9c",x"4c",x"70"),
   697 => (x"fb",x"c0",x"87",x"d8"),
   698 => (x"87",x"d2",x"02",x"ac"),
   699 => (x"d1",x"ef",x"55",x"74"),
   700 => (x"9c",x"4c",x"70",x"87"),
   701 => (x"c0",x"87",x"c7",x"02"),
   702 => (x"ff",x"05",x"ac",x"fb"),
   703 => (x"e0",x"c0",x"87",x"ee"),
   704 => (x"55",x"c1",x"c2",x"55"),
   705 => (x"d8",x"7d",x"97",x"c0"),
   706 => (x"a9",x"6e",x"49",x"66"),
   707 => (x"c8",x"87",x"db",x"05"),
   708 => (x"66",x"cc",x"48",x"66"),
   709 => (x"87",x"ca",x"04",x"a8"),
   710 => (x"c1",x"48",x"66",x"c8"),
   711 => (x"58",x"a6",x"cc",x"80"),
   712 => (x"66",x"cc",x"87",x"c8"),
   713 => (x"d0",x"88",x"c1",x"48"),
   714 => (x"d5",x"ee",x"58",x"a6"),
   715 => (x"c1",x"4c",x"70",x"87"),
   716 => (x"c8",x"05",x"ac",x"d0"),
   717 => (x"48",x"66",x"d4",x"87"),
   718 => (x"a6",x"d8",x"80",x"c1"),
   719 => (x"ac",x"d0",x"c1",x"58"),
   720 => (x"87",x"ea",x"fd",x"02"),
   721 => (x"48",x"a6",x"e0",x"c0"),
   722 => (x"c4",x"78",x"66",x"d8"),
   723 => (x"e0",x"c0",x"48",x"66"),
   724 => (x"c9",x"05",x"a8",x"66"),
   725 => (x"e4",x"c0",x"87",x"d8"),
   726 => (x"78",x"c0",x"48",x"a6"),
   727 => (x"78",x"c0",x"80",x"c4"),
   728 => (x"fb",x"c0",x"48",x"74"),
   729 => (x"6e",x"7e",x"70",x"88"),
   730 => (x"87",x"db",x"c8",x"02"),
   731 => (x"88",x"cb",x"48",x"6e"),
   732 => (x"02",x"6e",x"7e",x"70"),
   733 => (x"6e",x"87",x"ca",x"c1"),
   734 => (x"70",x"88",x"c9",x"48"),
   735 => (x"c3",x"02",x"6e",x"7e"),
   736 => (x"48",x"6e",x"87",x"e3"),
   737 => (x"7e",x"70",x"88",x"c4"),
   738 => (x"87",x"ce",x"02",x"6e"),
   739 => (x"88",x"c1",x"48",x"6e"),
   740 => (x"02",x"6e",x"7e",x"70"),
   741 => (x"c7",x"87",x"ce",x"c3"),
   742 => (x"a6",x"dc",x"87",x"e8"),
   743 => (x"78",x"f0",x"c0",x"48"),
   744 => (x"70",x"87",x"df",x"ec"),
   745 => (x"ac",x"ec",x"c0",x"4c"),
   746 => (x"c0",x"87",x"c4",x"02"),
   747 => (x"c0",x"5c",x"a6",x"e0"),
   748 => (x"cc",x"02",x"ac",x"ec"),
   749 => (x"87",x"ca",x"ec",x"87"),
   750 => (x"ec",x"c0",x"4c",x"70"),
   751 => (x"f4",x"ff",x"05",x"ac"),
   752 => (x"ac",x"ec",x"c0",x"87"),
   753 => (x"87",x"c3",x"c0",x"02"),
   754 => (x"c0",x"87",x"f7",x"eb"),
   755 => (x"d0",x"1e",x"ca",x"1e"),
   756 => (x"91",x"cb",x"49",x"66"),
   757 => (x"48",x"66",x"c8",x"c1"),
   758 => (x"a6",x"cc",x"80",x"71"),
   759 => (x"48",x"66",x"c8",x"58"),
   760 => (x"a6",x"d0",x"80",x"c4"),
   761 => (x"bf",x"66",x"cc",x"58"),
   762 => (x"87",x"da",x"ec",x"49"),
   763 => (x"1e",x"de",x"1e",x"c1"),
   764 => (x"49",x"bf",x"66",x"d4"),
   765 => (x"d0",x"87",x"cf",x"ec"),
   766 => (x"c0",x"49",x"70",x"86"),
   767 => (x"ec",x"c0",x"89",x"09"),
   768 => (x"e8",x"c0",x"59",x"a6"),
   769 => (x"a8",x"c0",x"48",x"66"),
   770 => (x"87",x"ee",x"c0",x"06"),
   771 => (x"48",x"66",x"e8",x"c0"),
   772 => (x"c0",x"03",x"a8",x"dd"),
   773 => (x"66",x"c4",x"87",x"e4"),
   774 => (x"e8",x"c0",x"49",x"bf"),
   775 => (x"e0",x"c0",x"81",x"66"),
   776 => (x"66",x"e8",x"c0",x"51"),
   777 => (x"c4",x"81",x"c1",x"49"),
   778 => (x"c2",x"81",x"bf",x"66"),
   779 => (x"e8",x"c0",x"51",x"c1"),
   780 => (x"81",x"c2",x"49",x"66"),
   781 => (x"81",x"bf",x"66",x"c4"),
   782 => (x"48",x"6e",x"51",x"c0"),
   783 => (x"78",x"cf",x"e2",x"c0"),
   784 => (x"81",x"c8",x"49",x"6e"),
   785 => (x"6e",x"51",x"66",x"d0"),
   786 => (x"d4",x"81",x"c9",x"49"),
   787 => (x"49",x"6e",x"51",x"66"),
   788 => (x"66",x"dc",x"81",x"ca"),
   789 => (x"48",x"66",x"d0",x"51"),
   790 => (x"a6",x"d4",x"80",x"c1"),
   791 => (x"80",x"d8",x"48",x"58"),
   792 => (x"e2",x"c4",x"78",x"c1"),
   793 => (x"87",x"cd",x"ec",x"87"),
   794 => (x"ec",x"c0",x"49",x"70"),
   795 => (x"c4",x"ec",x"59",x"a6"),
   796 => (x"c0",x"49",x"70",x"87"),
   797 => (x"dc",x"59",x"a6",x"e0"),
   798 => (x"ec",x"c0",x"48",x"66"),
   799 => (x"ca",x"c0",x"05",x"a8"),
   800 => (x"48",x"a6",x"dc",x"87"),
   801 => (x"78",x"66",x"e8",x"c0"),
   802 => (x"e8",x"87",x"c3",x"c0"),
   803 => (x"66",x"c8",x"87",x"f4"),
   804 => (x"c1",x"91",x"cb",x"49"),
   805 => (x"71",x"48",x"66",x"c0"),
   806 => (x"6e",x"7e",x"70",x"80"),
   807 => (x"6e",x"82",x"c8",x"4a"),
   808 => (x"c0",x"81",x"ca",x"49"),
   809 => (x"dc",x"51",x"66",x"e8"),
   810 => (x"81",x"c1",x"49",x"66"),
   811 => (x"89",x"66",x"e8",x"c0"),
   812 => (x"30",x"71",x"48",x"c1"),
   813 => (x"89",x"c1",x"49",x"70"),
   814 => (x"c1",x"7a",x"97",x"71"),
   815 => (x"49",x"bf",x"d6",x"fa"),
   816 => (x"29",x"66",x"e8",x"c0"),
   817 => (x"48",x"4a",x"6a",x"97"),
   818 => (x"f0",x"c0",x"98",x"71"),
   819 => (x"49",x"6e",x"58",x"a6"),
   820 => (x"4d",x"69",x"81",x"c4"),
   821 => (x"48",x"66",x"e0",x"c0"),
   822 => (x"02",x"a8",x"66",x"c4"),
   823 => (x"c4",x"87",x"c8",x"c0"),
   824 => (x"78",x"c0",x"48",x"a6"),
   825 => (x"c4",x"87",x"c5",x"c0"),
   826 => (x"78",x"c1",x"48",x"a6"),
   827 => (x"c0",x"1e",x"66",x"c4"),
   828 => (x"49",x"75",x"1e",x"e0"),
   829 => (x"c8",x"87",x"cf",x"e8"),
   830 => (x"c0",x"4c",x"70",x"86"),
   831 => (x"c1",x"06",x"ac",x"b7"),
   832 => (x"85",x"74",x"87",x"d3"),
   833 => (x"74",x"49",x"e0",x"c0"),
   834 => (x"c0",x"4b",x"75",x"89"),
   835 => (x"71",x"4a",x"db",x"f8"),
   836 => (x"87",x"d5",x"cd",x"ff"),
   837 => (x"e4",x"c0",x"85",x"c2"),
   838 => (x"80",x"c1",x"48",x"66"),
   839 => (x"58",x"a6",x"e8",x"c0"),
   840 => (x"49",x"66",x"ec",x"c0"),
   841 => (x"a9",x"70",x"81",x"c1"),
   842 => (x"87",x"c8",x"c0",x"02"),
   843 => (x"c0",x"48",x"a6",x"c4"),
   844 => (x"87",x"c5",x"c0",x"78"),
   845 => (x"c1",x"48",x"a6",x"c4"),
   846 => (x"1e",x"66",x"c4",x"78"),
   847 => (x"c0",x"49",x"a4",x"c2"),
   848 => (x"88",x"71",x"48",x"e0"),
   849 => (x"75",x"1e",x"49",x"70"),
   850 => (x"87",x"fa",x"e6",x"49"),
   851 => (x"b7",x"c0",x"86",x"c8"),
   852 => (x"c1",x"ff",x"01",x"a8"),
   853 => (x"66",x"e4",x"c0",x"87"),
   854 => (x"87",x"d1",x"c0",x"02"),
   855 => (x"81",x"c9",x"49",x"6e"),
   856 => (x"51",x"66",x"e4",x"c0"),
   857 => (x"e3",x"c0",x"48",x"6e"),
   858 => (x"cc",x"c0",x"78",x"e7"),
   859 => (x"c9",x"49",x"6e",x"87"),
   860 => (x"6e",x"51",x"c2",x"81"),
   861 => (x"db",x"e4",x"c0",x"48"),
   862 => (x"a6",x"e8",x"c0",x"78"),
   863 => (x"c0",x"78",x"c1",x"48"),
   864 => (x"ed",x"e5",x"87",x"c5"),
   865 => (x"c0",x"4c",x"70",x"87"),
   866 => (x"c0",x"02",x"66",x"e8"),
   867 => (x"66",x"c8",x"87",x"f4"),
   868 => (x"a8",x"66",x"cc",x"48"),
   869 => (x"87",x"cb",x"c0",x"04"),
   870 => (x"c1",x"48",x"66",x"c8"),
   871 => (x"58",x"a6",x"cc",x"80"),
   872 => (x"cc",x"87",x"df",x"c0"),
   873 => (x"88",x"c1",x"48",x"66"),
   874 => (x"c0",x"58",x"a6",x"d0"),
   875 => (x"c6",x"c1",x"87",x"d4"),
   876 => (x"c8",x"c0",x"05",x"ac"),
   877 => (x"48",x"66",x"d0",x"87"),
   878 => (x"a6",x"d4",x"80",x"c1"),
   879 => (x"87",x"f2",x"e4",x"58"),
   880 => (x"66",x"d4",x"4c",x"70"),
   881 => (x"d8",x"80",x"c1",x"48"),
   882 => (x"9c",x"74",x"58",x"a6"),
   883 => (x"87",x"cb",x"c0",x"02"),
   884 => (x"c1",x"48",x"66",x"c8"),
   885 => (x"04",x"a8",x"66",x"c8"),
   886 => (x"e4",x"87",x"fe",x"f2"),
   887 => (x"66",x"c8",x"87",x"cb"),
   888 => (x"03",x"a8",x"c7",x"48"),
   889 => (x"c1",x"87",x"e5",x"c0"),
   890 => (x"c0",x"48",x"f6",x"f6"),
   891 => (x"49",x"66",x"c8",x"78"),
   892 => (x"c0",x"c1",x"91",x"cb"),
   893 => (x"a1",x"c4",x"81",x"66"),
   894 => (x"c0",x"4a",x"6a",x"4a"),
   895 => (x"66",x"c8",x"79",x"52"),
   896 => (x"cc",x"80",x"c1",x"48"),
   897 => (x"a8",x"c7",x"58",x"a6"),
   898 => (x"87",x"db",x"ff",x"04"),
   899 => (x"e9",x"8e",x"d0",x"ff"),
   900 => (x"6f",x"4c",x"87",x"f5"),
   901 => (x"2a",x"20",x"64",x"61"),
   902 => (x"3a",x"00",x"20",x"2e"),
   903 => (x"73",x"1e",x"00",x"20"),
   904 => (x"9b",x"4b",x"71",x"1e"),
   905 => (x"c1",x"87",x"c6",x"02"),
   906 => (x"c0",x"48",x"f2",x"f6"),
   907 => (x"c1",x"1e",x"c7",x"78"),
   908 => (x"49",x"bf",x"f2",x"f6"),
   909 => (x"d6",x"fa",x"c0",x"1e"),
   910 => (x"ee",x"f6",x"c1",x"1e"),
   911 => (x"c0",x"ee",x"49",x"bf"),
   912 => (x"c1",x"86",x"cc",x"87"),
   913 => (x"49",x"bf",x"ee",x"f6"),
   914 => (x"73",x"87",x"f4",x"e9"),
   915 => (x"87",x"c8",x"02",x"9b"),
   916 => (x"49",x"d6",x"fa",x"c0"),
   917 => (x"87",x"e4",x"e2",x"c0"),
   918 => (x"1e",x"87",x"f0",x"e8"),
   919 => (x"c1",x"87",x"f1",x"c5"),
   920 => (x"87",x"fa",x"fe",x"49"),
   921 => (x"26",x"87",x"e8",x"c2"),
   922 => (x"e6",x"c0",x"1e",x"4f"),
   923 => (x"87",x"fa",x"87",x"ea"),
   924 => (x"c1",x"1e",x"4f",x"26"),
   925 => (x"c0",x"48",x"f2",x"f6"),
   926 => (x"ee",x"f6",x"c1",x"78"),
   927 => (x"ff",x"78",x"c0",x"48"),
   928 => (x"87",x"e5",x"87",x"d9"),
   929 => (x"4f",x"26",x"48",x"c0"),
   930 => (x"78",x"45",x"20",x"80"),
   931 => (x"80",x"00",x"74",x"69"),
   932 => (x"63",x"61",x"42",x"20"),
   933 => (x"08",x"97",x"00",x"6b"),
   934 => (x"1d",x"ba",x"00",x"00"),
   935 => (x"00",x"00",x"00",x"00"),
   936 => (x"00",x"08",x"97",x"00"),
   937 => (x"00",x"1d",x"d8",x"00"),
   938 => (x"00",x"00",x"00",x"00"),
   939 => (x"00",x"00",x"08",x"97"),
   940 => (x"00",x"00",x"1d",x"f6"),
   941 => (x"97",x"00",x"00",x"00"),
   942 => (x"14",x"00",x"00",x"08"),
   943 => (x"00",x"00",x"00",x"1e"),
   944 => (x"08",x"97",x"00",x"00"),
   945 => (x"1e",x"32",x"00",x"00"),
   946 => (x"00",x"00",x"00",x"00"),
   947 => (x"00",x"08",x"97",x"00"),
   948 => (x"00",x"1e",x"50",x"00"),
   949 => (x"00",x"00",x"00",x"00"),
   950 => (x"00",x"00",x"08",x"97"),
   951 => (x"00",x"00",x"1e",x"6e"),
   952 => (x"97",x"00",x"00",x"00"),
   953 => (x"00",x"00",x"00",x"08"),
   954 => (x"00",x"00",x"00",x"00"),
   955 => (x"09",x"32",x"00",x"00"),
   956 => (x"00",x"00",x"00",x"00"),
   957 => (x"00",x"00",x"00",x"00"),
   958 => (x"f0",x"fe",x"1e",x"00"),
   959 => (x"cd",x"78",x"c0",x"48"),
   960 => (x"26",x"09",x"79",x"09"),
   961 => (x"fe",x"1e",x"1e",x"4f"),
   962 => (x"48",x"7e",x"bf",x"f0"),
   963 => (x"1e",x"4f",x"26",x"26"),
   964 => (x"c1",x"48",x"f0",x"fe"),
   965 => (x"1e",x"4f",x"26",x"78"),
   966 => (x"c0",x"48",x"f0",x"fe"),
   967 => (x"1e",x"4f",x"26",x"78"),
   968 => (x"52",x"c0",x"4a",x"71"),
   969 => (x"0e",x"4f",x"26",x"52"),
   970 => (x"5d",x"5c",x"5b",x"5e"),
   971 => (x"71",x"86",x"f4",x"0e"),
   972 => (x"7e",x"6d",x"97",x"4d"),
   973 => (x"97",x"4c",x"a5",x"c1"),
   974 => (x"a6",x"c8",x"48",x"6c"),
   975 => (x"c4",x"48",x"6e",x"58"),
   976 => (x"c5",x"05",x"a8",x"66"),
   977 => (x"c0",x"48",x"ff",x"87"),
   978 => (x"ca",x"ff",x"87",x"e6"),
   979 => (x"49",x"a5",x"c2",x"87"),
   980 => (x"71",x"4b",x"6c",x"97"),
   981 => (x"6b",x"97",x"4b",x"a3"),
   982 => (x"7e",x"6c",x"97",x"4b"),
   983 => (x"80",x"c1",x"48",x"6e"),
   984 => (x"c7",x"58",x"a6",x"c8"),
   985 => (x"58",x"a6",x"cc",x"98"),
   986 => (x"fe",x"7c",x"97",x"70"),
   987 => (x"48",x"73",x"87",x"e1"),
   988 => (x"4d",x"26",x"8e",x"f4"),
   989 => (x"4b",x"26",x"4c",x"26"),
   990 => (x"5e",x"0e",x"4f",x"26"),
   991 => (x"f4",x"0e",x"5c",x"5b"),
   992 => (x"d8",x"4c",x"71",x"86"),
   993 => (x"ff",x"c3",x"4a",x"66"),
   994 => (x"4b",x"a4",x"c2",x"9a"),
   995 => (x"73",x"49",x"6c",x"97"),
   996 => (x"51",x"72",x"49",x"a1"),
   997 => (x"6e",x"7e",x"6c",x"97"),
   998 => (x"c8",x"80",x"c1",x"48"),
   999 => (x"98",x"c7",x"58",x"a6"),
  1000 => (x"70",x"58",x"a6",x"cc"),
  1001 => (x"ff",x"8e",x"f4",x"54"),
  1002 => (x"1e",x"1e",x"87",x"ca"),
  1003 => (x"e0",x"87",x"e8",x"fd"),
  1004 => (x"c0",x"49",x"4a",x"bf"),
  1005 => (x"02",x"99",x"c0",x"e0"),
  1006 => (x"1e",x"72",x"87",x"cb"),
  1007 => (x"49",x"cc",x"fa",x"c1"),
  1008 => (x"c4",x"87",x"f7",x"fe"),
  1009 => (x"87",x"fd",x"fc",x"86"),
  1010 => (x"c2",x"fd",x"7e",x"70"),
  1011 => (x"4f",x"26",x"26",x"87"),
  1012 => (x"cc",x"fa",x"c1",x"1e"),
  1013 => (x"87",x"c7",x"fd",x"49"),
  1014 => (x"49",x"ea",x"fe",x"c0"),
  1015 => (x"c4",x"87",x"da",x"fc"),
  1016 => (x"4f",x"26",x"87",x"c1"),
  1017 => (x"48",x"d0",x"ff",x"1e"),
  1018 => (x"ff",x"78",x"e1",x"c8"),
  1019 => (x"78",x"c5",x"48",x"d4"),
  1020 => (x"bf",x"f6",x"c5",x"c1"),
  1021 => (x"c3",x"87",x"c3",x"02"),
  1022 => (x"66",x"c8",x"78",x"e0"),
  1023 => (x"ff",x"87",x"c6",x"02"),
  1024 => (x"f0",x"c3",x"48",x"d4"),
  1025 => (x"48",x"d4",x"ff",x"78"),
  1026 => (x"d0",x"ff",x"78",x"71"),
  1027 => (x"78",x"e1",x"c8",x"48"),
  1028 => (x"26",x"78",x"e0",x"c0"),
  1029 => (x"5b",x"5e",x"0e",x"4f"),
  1030 => (x"4c",x"71",x"0e",x"5c"),
  1031 => (x"49",x"cc",x"fa",x"c1"),
  1032 => (x"70",x"87",x"c4",x"fc"),
  1033 => (x"aa",x"b7",x"c0",x"4a"),
  1034 => (x"87",x"e2",x"c2",x"04"),
  1035 => (x"05",x"aa",x"f0",x"c3"),
  1036 => (x"c5",x"c1",x"87",x"c9"),
  1037 => (x"78",x"c1",x"48",x"f2"),
  1038 => (x"c3",x"87",x"c3",x"c2"),
  1039 => (x"c9",x"05",x"aa",x"e0"),
  1040 => (x"f6",x"c5",x"c1",x"87"),
  1041 => (x"c1",x"78",x"c1",x"48"),
  1042 => (x"c5",x"c1",x"87",x"f4"),
  1043 => (x"c6",x"02",x"bf",x"f6"),
  1044 => (x"a2",x"c0",x"c2",x"87"),
  1045 => (x"72",x"87",x"c2",x"4b"),
  1046 => (x"05",x"9c",x"74",x"4b"),
  1047 => (x"c5",x"c1",x"87",x"d1"),
  1048 => (x"c1",x"1e",x"bf",x"f2"),
  1049 => (x"1e",x"bf",x"f6",x"c5"),
  1050 => (x"f7",x"fd",x"49",x"72"),
  1051 => (x"c1",x"86",x"c8",x"87"),
  1052 => (x"02",x"bf",x"f2",x"c5"),
  1053 => (x"73",x"87",x"e0",x"c0"),
  1054 => (x"29",x"b7",x"c4",x"49"),
  1055 => (x"f2",x"c4",x"c1",x"91"),
  1056 => (x"cf",x"4a",x"73",x"81"),
  1057 => (x"c1",x"92",x"c2",x"9a"),
  1058 => (x"70",x"30",x"72",x"48"),
  1059 => (x"72",x"ba",x"ff",x"4a"),
  1060 => (x"70",x"98",x"69",x"48"),
  1061 => (x"73",x"87",x"db",x"79"),
  1062 => (x"29",x"b7",x"c4",x"49"),
  1063 => (x"f2",x"c4",x"c1",x"91"),
  1064 => (x"cf",x"4a",x"73",x"81"),
  1065 => (x"c3",x"92",x"c2",x"9a"),
  1066 => (x"70",x"30",x"72",x"48"),
  1067 => (x"b0",x"69",x"48",x"4a"),
  1068 => (x"c5",x"c1",x"79",x"70"),
  1069 => (x"78",x"c0",x"48",x"f6"),
  1070 => (x"48",x"f2",x"c5",x"c1"),
  1071 => (x"fa",x"c1",x"78",x"c0"),
  1072 => (x"e2",x"f9",x"49",x"cc"),
  1073 => (x"c0",x"4a",x"70",x"87"),
  1074 => (x"fd",x"03",x"aa",x"b7"),
  1075 => (x"48",x"c0",x"87",x"de"),
  1076 => (x"4d",x"26",x"87",x"c2"),
  1077 => (x"4b",x"26",x"4c",x"26"),
  1078 => (x"71",x"1e",x"4f",x"26"),
  1079 => (x"f4",x"fc",x"49",x"4a"),
  1080 => (x"1e",x"4f",x"26",x"87"),
  1081 => (x"49",x"72",x"4a",x"c0"),
  1082 => (x"c4",x"c1",x"91",x"c4"),
  1083 => (x"79",x"c0",x"81",x"f2"),
  1084 => (x"b7",x"d0",x"82",x"c1"),
  1085 => (x"87",x"ee",x"04",x"aa"),
  1086 => (x"5e",x"0e",x"4f",x"26"),
  1087 => (x"0e",x"5d",x"5c",x"5b"),
  1088 => (x"d2",x"f8",x"4d",x"71"),
  1089 => (x"c4",x"4a",x"75",x"87"),
  1090 => (x"c1",x"92",x"2a",x"b7"),
  1091 => (x"75",x"82",x"f2",x"c4"),
  1092 => (x"c2",x"9c",x"cf",x"4c"),
  1093 => (x"4b",x"49",x"6a",x"94"),
  1094 => (x"9b",x"c3",x"2b",x"74"),
  1095 => (x"30",x"74",x"48",x"c2"),
  1096 => (x"bc",x"ff",x"4c",x"70"),
  1097 => (x"98",x"71",x"48",x"74"),
  1098 => (x"e2",x"f7",x"7a",x"70"),
  1099 => (x"fe",x"48",x"73",x"87"),
  1100 => (x"00",x"00",x"87",x"e0"),
  1101 => (x"30",x"30",x"00",x"00"),
  1102 => (x"30",x"30",x"30",x"30"),
  1103 => (x"30",x"30",x"30",x"30"),
  1104 => (x"30",x"30",x"30",x"30"),
  1105 => (x"30",x"30",x"30",x"30"),
  1106 => (x"30",x"30",x"30",x"30"),
  1107 => (x"30",x"30",x"30",x"30"),
  1108 => (x"30",x"30",x"30",x"30"),
  1109 => (x"30",x"30",x"30",x"30"),
  1110 => (x"30",x"30",x"30",x"30"),
  1111 => (x"30",x"30",x"30",x"30"),
  1112 => (x"30",x"30",x"30",x"30"),
  1113 => (x"30",x"30",x"30",x"30"),
  1114 => (x"30",x"30",x"30",x"30"),
  1115 => (x"30",x"30",x"30",x"30"),
  1116 => (x"00",x"00",x"30",x"30"),
  1117 => (x"00",x"00",x"00",x"00"),
  1118 => (x"ff",x"1e",x"00",x"00"),
  1119 => (x"e1",x"c8",x"48",x"d0"),
  1120 => (x"ff",x"48",x"71",x"78"),
  1121 => (x"c4",x"78",x"08",x"d4"),
  1122 => (x"d4",x"ff",x"48",x"66"),
  1123 => (x"4f",x"26",x"78",x"08"),
  1124 => (x"c4",x"4a",x"71",x"1e"),
  1125 => (x"72",x"1e",x"49",x"66"),
  1126 => (x"87",x"de",x"ff",x"49"),
  1127 => (x"c0",x"48",x"d0",x"ff"),
  1128 => (x"26",x"26",x"78",x"e0"),
  1129 => (x"1e",x"73",x"1e",x"4f"),
  1130 => (x"66",x"c8",x"4b",x"71"),
  1131 => (x"4a",x"73",x"1e",x"49"),
  1132 => (x"49",x"a2",x"e0",x"c1"),
  1133 => (x"26",x"87",x"d9",x"ff"),
  1134 => (x"4d",x"26",x"87",x"c4"),
  1135 => (x"4b",x"26",x"4c",x"26"),
  1136 => (x"73",x"1e",x"4f",x"26"),
  1137 => (x"4b",x"4a",x"71",x"1e"),
  1138 => (x"03",x"ab",x"b7",x"c2"),
  1139 => (x"49",x"a3",x"87",x"c8"),
  1140 => (x"9a",x"ff",x"c3",x"4a"),
  1141 => (x"a3",x"ce",x"87",x"c7"),
  1142 => (x"ff",x"c3",x"4a",x"49"),
  1143 => (x"49",x"66",x"c8",x"9a"),
  1144 => (x"fe",x"49",x"72",x"1e"),
  1145 => (x"ff",x"26",x"87",x"ea"),
  1146 => (x"ff",x"1e",x"87",x"d4"),
  1147 => (x"ff",x"c3",x"4a",x"d4"),
  1148 => (x"48",x"d0",x"ff",x"7a"),
  1149 => (x"de",x"78",x"e1",x"c0"),
  1150 => (x"d6",x"fa",x"c1",x"7a"),
  1151 => (x"48",x"49",x"7a",x"bf"),
  1152 => (x"7a",x"70",x"28",x"c8"),
  1153 => (x"28",x"d0",x"48",x"71"),
  1154 => (x"48",x"71",x"7a",x"70"),
  1155 => (x"7a",x"70",x"28",x"d8"),
  1156 => (x"c0",x"48",x"d0",x"ff"),
  1157 => (x"4f",x"26",x"78",x"e0"),
  1158 => (x"5c",x"5b",x"5e",x"0e"),
  1159 => (x"4c",x"71",x"0e",x"5d"),
  1160 => (x"bf",x"d6",x"fa",x"c1"),
  1161 => (x"2b",x"74",x"4b",x"4d"),
  1162 => (x"c1",x"9b",x"66",x"d0"),
  1163 => (x"ab",x"66",x"d4",x"83"),
  1164 => (x"c0",x"87",x"c2",x"04"),
  1165 => (x"d0",x"4a",x"74",x"4b"),
  1166 => (x"31",x"72",x"49",x"66"),
  1167 => (x"99",x"75",x"b9",x"ff"),
  1168 => (x"30",x"72",x"48",x"73"),
  1169 => (x"71",x"48",x"4a",x"70"),
  1170 => (x"da",x"fa",x"c1",x"b0"),
  1171 => (x"87",x"da",x"fe",x"58"),
  1172 => (x"4c",x"26",x"4d",x"26"),
  1173 => (x"4f",x"26",x"4b",x"26"),
  1174 => (x"48",x"d0",x"ff",x"1e"),
  1175 => (x"71",x"78",x"c9",x"c8"),
  1176 => (x"08",x"d4",x"ff",x"48"),
  1177 => (x"1e",x"4f",x"26",x"78"),
  1178 => (x"eb",x"49",x"4a",x"71"),
  1179 => (x"48",x"d0",x"ff",x"87"),
  1180 => (x"4f",x"26",x"78",x"c8"),
  1181 => (x"71",x"1e",x"73",x"1e"),
  1182 => (x"e6",x"fa",x"c1",x"4b"),
  1183 => (x"87",x"c3",x"02",x"bf"),
  1184 => (x"ff",x"87",x"eb",x"c2"),
  1185 => (x"c9",x"c8",x"48",x"d0"),
  1186 => (x"c0",x"49",x"73",x"78"),
  1187 => (x"d4",x"ff",x"b1",x"e0"),
  1188 => (x"c1",x"78",x"71",x"48"),
  1189 => (x"c0",x"48",x"da",x"fa"),
  1190 => (x"02",x"66",x"c8",x"78"),
  1191 => (x"ff",x"c3",x"87",x"c5"),
  1192 => (x"c0",x"87",x"c2",x"49"),
  1193 => (x"e2",x"fa",x"c1",x"49"),
  1194 => (x"02",x"66",x"cc",x"59"),
  1195 => (x"d5",x"c5",x"87",x"c6"),
  1196 => (x"87",x"c4",x"4a",x"d5"),
  1197 => (x"4a",x"ff",x"ff",x"cf"),
  1198 => (x"5a",x"e6",x"fa",x"c1"),
  1199 => (x"48",x"e6",x"fa",x"c1"),
  1200 => (x"87",x"c4",x"78",x"c1"),
  1201 => (x"4c",x"26",x"4d",x"26"),
  1202 => (x"4f",x"26",x"4b",x"26"),
  1203 => (x"5c",x"5b",x"5e",x"0e"),
  1204 => (x"4a",x"71",x"0e",x"5d"),
  1205 => (x"bf",x"e2",x"fa",x"c1"),
  1206 => (x"02",x"9a",x"72",x"4c"),
  1207 => (x"c8",x"49",x"87",x"cb"),
  1208 => (x"ea",x"c9",x"c1",x"91"),
  1209 => (x"c4",x"83",x"71",x"4b"),
  1210 => (x"ea",x"cd",x"c1",x"87"),
  1211 => (x"13",x"4d",x"c0",x"4b"),
  1212 => (x"c1",x"99",x"74",x"49"),
  1213 => (x"b9",x"bf",x"de",x"fa"),
  1214 => (x"71",x"48",x"d4",x"ff"),
  1215 => (x"2c",x"b7",x"c1",x"78"),
  1216 => (x"ad",x"b7",x"c8",x"85"),
  1217 => (x"c1",x"87",x"e8",x"04"),
  1218 => (x"48",x"bf",x"da",x"fa"),
  1219 => (x"fa",x"c1",x"80",x"c8"),
  1220 => (x"ef",x"fe",x"58",x"de"),
  1221 => (x"1e",x"73",x"1e",x"87"),
  1222 => (x"4a",x"13",x"4b",x"71"),
  1223 => (x"87",x"cb",x"02",x"9a"),
  1224 => (x"e7",x"fe",x"49",x"72"),
  1225 => (x"9a",x"4a",x"13",x"87"),
  1226 => (x"fe",x"87",x"f5",x"05"),
  1227 => (x"c1",x"1e",x"87",x"da"),
  1228 => (x"49",x"bf",x"da",x"fa"),
  1229 => (x"48",x"da",x"fa",x"c1"),
  1230 => (x"c4",x"78",x"a1",x"c1"),
  1231 => (x"03",x"a9",x"b7",x"c0"),
  1232 => (x"d4",x"ff",x"87",x"db"),
  1233 => (x"de",x"fa",x"c1",x"48"),
  1234 => (x"fa",x"c1",x"78",x"bf"),
  1235 => (x"c1",x"49",x"bf",x"da"),
  1236 => (x"c1",x"48",x"da",x"fa"),
  1237 => (x"c0",x"c4",x"78",x"a1"),
  1238 => (x"e5",x"04",x"a9",x"b7"),
  1239 => (x"48",x"d0",x"ff",x"87"),
  1240 => (x"fa",x"c1",x"78",x"c8"),
  1241 => (x"78",x"c0",x"48",x"e6"),
  1242 => (x"00",x"00",x"4f",x"26"),
  1243 => (x"00",x"00",x"00",x"00"),
  1244 => (x"00",x"00",x"00",x"00"),
  1245 => (x"00",x"5f",x"5f",x"00"),
  1246 => (x"03",x"00",x"00",x"00"),
  1247 => (x"03",x"03",x"00",x"03"),
  1248 => (x"7f",x"14",x"00",x"00"),
  1249 => (x"7f",x"7f",x"14",x"7f"),
  1250 => (x"24",x"00",x"00",x"14"),
  1251 => (x"3a",x"6b",x"6b",x"2e"),
  1252 => (x"6a",x"4c",x"00",x"12"),
  1253 => (x"56",x"6c",x"18",x"36"),
  1254 => (x"7e",x"30",x"00",x"32"),
  1255 => (x"3a",x"77",x"59",x"4f"),
  1256 => (x"00",x"00",x"40",x"68"),
  1257 => (x"00",x"03",x"07",x"04"),
  1258 => (x"00",x"00",x"00",x"00"),
  1259 => (x"41",x"63",x"3e",x"1c"),
  1260 => (x"00",x"00",x"00",x"00"),
  1261 => (x"1c",x"3e",x"63",x"41"),
  1262 => (x"2a",x"08",x"00",x"00"),
  1263 => (x"3e",x"1c",x"1c",x"3e"),
  1264 => (x"08",x"00",x"08",x"2a"),
  1265 => (x"08",x"3e",x"3e",x"08"),
  1266 => (x"00",x"00",x"00",x"08"),
  1267 => (x"00",x"60",x"e0",x"80"),
  1268 => (x"08",x"00",x"00",x"00"),
  1269 => (x"08",x"08",x"08",x"08"),
  1270 => (x"00",x"00",x"00",x"08"),
  1271 => (x"00",x"60",x"60",x"00"),
  1272 => (x"60",x"40",x"00",x"00"),
  1273 => (x"06",x"0c",x"18",x"30"),
  1274 => (x"3e",x"00",x"01",x"03"),
  1275 => (x"7f",x"4d",x"59",x"7f"),
  1276 => (x"04",x"00",x"00",x"3e"),
  1277 => (x"00",x"7f",x"7f",x"06"),
  1278 => (x"42",x"00",x"00",x"00"),
  1279 => (x"4f",x"59",x"71",x"63"),
  1280 => (x"22",x"00",x"00",x"46"),
  1281 => (x"7f",x"49",x"49",x"63"),
  1282 => (x"1c",x"18",x"00",x"36"),
  1283 => (x"7f",x"7f",x"13",x"16"),
  1284 => (x"27",x"00",x"00",x"10"),
  1285 => (x"7d",x"45",x"45",x"67"),
  1286 => (x"3c",x"00",x"00",x"39"),
  1287 => (x"79",x"49",x"4b",x"7e"),
  1288 => (x"01",x"00",x"00",x"30"),
  1289 => (x"0f",x"79",x"71",x"01"),
  1290 => (x"36",x"00",x"00",x"07"),
  1291 => (x"7f",x"49",x"49",x"7f"),
  1292 => (x"06",x"00",x"00",x"36"),
  1293 => (x"3f",x"69",x"49",x"4f"),
  1294 => (x"00",x"00",x"00",x"1e"),
  1295 => (x"00",x"66",x"66",x"00"),
  1296 => (x"00",x"00",x"00",x"00"),
  1297 => (x"00",x"66",x"e6",x"80"),
  1298 => (x"08",x"00",x"00",x"00"),
  1299 => (x"22",x"14",x"14",x"08"),
  1300 => (x"14",x"00",x"00",x"22"),
  1301 => (x"14",x"14",x"14",x"14"),
  1302 => (x"22",x"00",x"00",x"14"),
  1303 => (x"08",x"14",x"14",x"22"),
  1304 => (x"02",x"00",x"00",x"08"),
  1305 => (x"0f",x"59",x"51",x"03"),
  1306 => (x"7f",x"3e",x"00",x"06"),
  1307 => (x"1f",x"55",x"5d",x"41"),
  1308 => (x"7e",x"00",x"00",x"1e"),
  1309 => (x"7f",x"09",x"09",x"7f"),
  1310 => (x"7f",x"00",x"00",x"7e"),
  1311 => (x"7f",x"49",x"49",x"7f"),
  1312 => (x"1c",x"00",x"00",x"36"),
  1313 => (x"41",x"41",x"63",x"3e"),
  1314 => (x"7f",x"00",x"00",x"41"),
  1315 => (x"3e",x"63",x"41",x"7f"),
  1316 => (x"7f",x"00",x"00",x"1c"),
  1317 => (x"41",x"49",x"49",x"7f"),
  1318 => (x"7f",x"00",x"00",x"41"),
  1319 => (x"01",x"09",x"09",x"7f"),
  1320 => (x"3e",x"00",x"00",x"01"),
  1321 => (x"7b",x"49",x"41",x"7f"),
  1322 => (x"7f",x"00",x"00",x"7a"),
  1323 => (x"7f",x"08",x"08",x"7f"),
  1324 => (x"00",x"00",x"00",x"7f"),
  1325 => (x"41",x"7f",x"7f",x"41"),
  1326 => (x"20",x"00",x"00",x"00"),
  1327 => (x"7f",x"40",x"40",x"60"),
  1328 => (x"7f",x"7f",x"00",x"3f"),
  1329 => (x"63",x"36",x"1c",x"08"),
  1330 => (x"7f",x"00",x"00",x"41"),
  1331 => (x"40",x"40",x"40",x"7f"),
  1332 => (x"7f",x"7f",x"00",x"40"),
  1333 => (x"7f",x"06",x"0c",x"06"),
  1334 => (x"7f",x"7f",x"00",x"7f"),
  1335 => (x"7f",x"18",x"0c",x"06"),
  1336 => (x"3e",x"00",x"00",x"7f"),
  1337 => (x"7f",x"41",x"41",x"7f"),
  1338 => (x"7f",x"00",x"00",x"3e"),
  1339 => (x"0f",x"09",x"09",x"7f"),
  1340 => (x"7f",x"3e",x"00",x"06"),
  1341 => (x"7e",x"7f",x"61",x"41"),
  1342 => (x"7f",x"00",x"00",x"40"),
  1343 => (x"7f",x"19",x"09",x"7f"),
  1344 => (x"26",x"00",x"00",x"66"),
  1345 => (x"7b",x"59",x"4d",x"6f"),
  1346 => (x"01",x"00",x"00",x"32"),
  1347 => (x"01",x"7f",x"7f",x"01"),
  1348 => (x"3f",x"00",x"00",x"01"),
  1349 => (x"7f",x"40",x"40",x"7f"),
  1350 => (x"0f",x"00",x"00",x"3f"),
  1351 => (x"3f",x"70",x"70",x"3f"),
  1352 => (x"7f",x"7f",x"00",x"0f"),
  1353 => (x"7f",x"30",x"18",x"30"),
  1354 => (x"63",x"41",x"00",x"7f"),
  1355 => (x"36",x"1c",x"1c",x"36"),
  1356 => (x"03",x"01",x"41",x"63"),
  1357 => (x"06",x"7c",x"7c",x"06"),
  1358 => (x"71",x"61",x"01",x"03"),
  1359 => (x"43",x"47",x"4d",x"59"),
  1360 => (x"00",x"00",x"00",x"41"),
  1361 => (x"41",x"41",x"7f",x"7f"),
  1362 => (x"03",x"01",x"00",x"00"),
  1363 => (x"30",x"18",x"0c",x"06"),
  1364 => (x"00",x"00",x"40",x"60"),
  1365 => (x"7f",x"7f",x"41",x"41"),
  1366 => (x"0c",x"08",x"00",x"00"),
  1367 => (x"0c",x"06",x"03",x"06"),
  1368 => (x"80",x"80",x"00",x"08"),
  1369 => (x"80",x"80",x"80",x"80"),
  1370 => (x"00",x"00",x"00",x"80"),
  1371 => (x"04",x"07",x"03",x"00"),
  1372 => (x"20",x"00",x"00",x"00"),
  1373 => (x"7c",x"54",x"54",x"74"),
  1374 => (x"7f",x"00",x"00",x"78"),
  1375 => (x"7c",x"44",x"44",x"7f"),
  1376 => (x"38",x"00",x"00",x"38"),
  1377 => (x"44",x"44",x"44",x"7c"),
  1378 => (x"38",x"00",x"00",x"00"),
  1379 => (x"7f",x"44",x"44",x"7c"),
  1380 => (x"38",x"00",x"00",x"7f"),
  1381 => (x"5c",x"54",x"54",x"7c"),
  1382 => (x"04",x"00",x"00",x"18"),
  1383 => (x"05",x"05",x"7f",x"7e"),
  1384 => (x"18",x"00",x"00",x"00"),
  1385 => (x"fc",x"a4",x"a4",x"bc"),
  1386 => (x"7f",x"00",x"00",x"7c"),
  1387 => (x"7c",x"04",x"04",x"7f"),
  1388 => (x"00",x"00",x"00",x"78"),
  1389 => (x"40",x"7d",x"3d",x"00"),
  1390 => (x"80",x"00",x"00",x"00"),
  1391 => (x"7d",x"fd",x"80",x"80"),
  1392 => (x"7f",x"00",x"00",x"00"),
  1393 => (x"6c",x"38",x"10",x"7f"),
  1394 => (x"00",x"00",x"00",x"44"),
  1395 => (x"40",x"7f",x"3f",x"00"),
  1396 => (x"7c",x"7c",x"00",x"00"),
  1397 => (x"7c",x"0c",x"18",x"0c"),
  1398 => (x"7c",x"00",x"00",x"78"),
  1399 => (x"7c",x"04",x"04",x"7c"),
  1400 => (x"38",x"00",x"00",x"78"),
  1401 => (x"7c",x"44",x"44",x"7c"),
  1402 => (x"fc",x"00",x"00",x"38"),
  1403 => (x"3c",x"24",x"24",x"fc"),
  1404 => (x"18",x"00",x"00",x"18"),
  1405 => (x"fc",x"24",x"24",x"3c"),
  1406 => (x"7c",x"00",x"00",x"fc"),
  1407 => (x"0c",x"04",x"04",x"7c"),
  1408 => (x"48",x"00",x"00",x"08"),
  1409 => (x"74",x"54",x"54",x"5c"),
  1410 => (x"04",x"00",x"00",x"20"),
  1411 => (x"44",x"44",x"7f",x"3f"),
  1412 => (x"3c",x"00",x"00",x"00"),
  1413 => (x"7c",x"40",x"40",x"7c"),
  1414 => (x"1c",x"00",x"00",x"7c"),
  1415 => (x"3c",x"60",x"60",x"3c"),
  1416 => (x"7c",x"3c",x"00",x"1c"),
  1417 => (x"7c",x"60",x"30",x"60"),
  1418 => (x"6c",x"44",x"00",x"3c"),
  1419 => (x"6c",x"38",x"10",x"38"),
  1420 => (x"1c",x"00",x"00",x"44"),
  1421 => (x"3c",x"60",x"e0",x"bc"),
  1422 => (x"44",x"00",x"00",x"1c"),
  1423 => (x"4c",x"5c",x"74",x"64"),
  1424 => (x"08",x"00",x"00",x"44"),
  1425 => (x"41",x"77",x"3e",x"08"),
  1426 => (x"00",x"00",x"00",x"41"),
  1427 => (x"00",x"7f",x"7f",x"00"),
  1428 => (x"41",x"00",x"00",x"00"),
  1429 => (x"08",x"3e",x"77",x"41"),
  1430 => (x"01",x"02",x"00",x"08"),
  1431 => (x"02",x"02",x"03",x"01"),
  1432 => (x"7f",x"7f",x"00",x"01"),
  1433 => (x"7f",x"7f",x"7f",x"7f"),
  1434 => (x"08",x"08",x"00",x"7f"),
  1435 => (x"3e",x"3e",x"1c",x"1c"),
  1436 => (x"7f",x"7f",x"7f",x"7f"),
  1437 => (x"1c",x"1c",x"3e",x"3e"),
  1438 => (x"10",x"00",x"08",x"08"),
  1439 => (x"18",x"7c",x"7c",x"18"),
  1440 => (x"10",x"00",x"00",x"10"),
  1441 => (x"30",x"7c",x"7c",x"30"),
  1442 => (x"30",x"10",x"00",x"10"),
  1443 => (x"1e",x"78",x"60",x"60"),
  1444 => (x"66",x"42",x"00",x"06"),
  1445 => (x"66",x"3c",x"18",x"3c"),
  1446 => (x"38",x"78",x"00",x"42"),
  1447 => (x"6c",x"c6",x"c2",x"6a"),
  1448 => (x"00",x"60",x"00",x"38"),
  1449 => (x"00",x"00",x"60",x"00"),
  1450 => (x"5e",x"0e",x"00",x"60"),
  1451 => (x"0e",x"5d",x"5c",x"5b"),
  1452 => (x"c1",x"4c",x"71",x"1e"),
  1453 => (x"4d",x"bf",x"f7",x"fa"),
  1454 => (x"1e",x"c0",x"4b",x"c0"),
  1455 => (x"c7",x"02",x"ab",x"74"),
  1456 => (x"48",x"a6",x"c4",x"87"),
  1457 => (x"87",x"c5",x"78",x"c0"),
  1458 => (x"c1",x"48",x"a6",x"c4"),
  1459 => (x"1e",x"66",x"c4",x"78"),
  1460 => (x"df",x"ee",x"49",x"73"),
  1461 => (x"c0",x"86",x"c8",x"87"),
  1462 => (x"ef",x"ef",x"49",x"e0"),
  1463 => (x"4a",x"a5",x"c4",x"87"),
  1464 => (x"f0",x"f0",x"49",x"6a"),
  1465 => (x"87",x"c6",x"f1",x"87"),
  1466 => (x"83",x"c1",x"85",x"cb"),
  1467 => (x"04",x"ab",x"b7",x"c8"),
  1468 => (x"26",x"87",x"c7",x"ff"),
  1469 => (x"4c",x"26",x"4d",x"26"),
  1470 => (x"4f",x"26",x"4b",x"26"),
  1471 => (x"c1",x"4a",x"71",x"1e"),
  1472 => (x"c1",x"5a",x"fb",x"fa"),
  1473 => (x"c7",x"48",x"fb",x"fa"),
  1474 => (x"dd",x"fe",x"49",x"78"),
  1475 => (x"1e",x"4f",x"26",x"87"),
  1476 => (x"4a",x"71",x"1e",x"73"),
  1477 => (x"03",x"aa",x"b7",x"c0"),
  1478 => (x"e8",x"c1",x"87",x"d3"),
  1479 => (x"c4",x"05",x"bf",x"cf"),
  1480 => (x"c2",x"4b",x"c1",x"87"),
  1481 => (x"c1",x"4b",x"c0",x"87"),
  1482 => (x"c4",x"5b",x"d3",x"e8"),
  1483 => (x"d3",x"e8",x"c1",x"87"),
  1484 => (x"cf",x"e8",x"c1",x"5a"),
  1485 => (x"9a",x"c1",x"4a",x"bf"),
  1486 => (x"49",x"a2",x"c0",x"c1"),
  1487 => (x"fc",x"87",x"e8",x"ec"),
  1488 => (x"cf",x"e8",x"c1",x"48"),
  1489 => (x"ef",x"fe",x"78",x"bf"),
  1490 => (x"4a",x"71",x"1e",x"87"),
  1491 => (x"72",x"1e",x"66",x"c4"),
  1492 => (x"87",x"ee",x"e9",x"49"),
  1493 => (x"1e",x"4f",x"26",x"26"),
  1494 => (x"bf",x"cf",x"e8",x"c1"),
  1495 => (x"87",x"fa",x"e5",x"49"),
  1496 => (x"48",x"ef",x"fa",x"c1"),
  1497 => (x"c1",x"78",x"bf",x"e8"),
  1498 => (x"ec",x"48",x"eb",x"fa"),
  1499 => (x"fa",x"c1",x"78",x"bf"),
  1500 => (x"49",x"4a",x"bf",x"ef"),
  1501 => (x"c8",x"99",x"ff",x"c3"),
  1502 => (x"48",x"72",x"2a",x"b7"),
  1503 => (x"fa",x"c1",x"b0",x"71"),
  1504 => (x"4f",x"26",x"58",x"f7"),
  1505 => (x"5c",x"5b",x"5e",x"0e"),
  1506 => (x"4b",x"71",x"0e",x"5d"),
  1507 => (x"c1",x"87",x"c8",x"ff"),
  1508 => (x"c0",x"48",x"ea",x"fa"),
  1509 => (x"e5",x"49",x"73",x"50"),
  1510 => (x"49",x"70",x"87",x"e0"),
  1511 => (x"cb",x"9c",x"c2",x"4c"),
  1512 => (x"f2",x"c9",x"49",x"ee"),
  1513 => (x"4d",x"49",x"70",x"87"),
  1514 => (x"97",x"ea",x"fa",x"c1"),
  1515 => (x"e2",x"c1",x"05",x"bf"),
  1516 => (x"49",x"66",x"d0",x"87"),
  1517 => (x"bf",x"f3",x"fa",x"c1"),
  1518 => (x"87",x"d6",x"05",x"99"),
  1519 => (x"c1",x"49",x"66",x"d4"),
  1520 => (x"99",x"bf",x"eb",x"fa"),
  1521 => (x"73",x"87",x"cb",x"05"),
  1522 => (x"87",x"ee",x"e4",x"49"),
  1523 => (x"c1",x"02",x"98",x"70"),
  1524 => (x"4c",x"c1",x"87",x"c1"),
  1525 => (x"75",x"87",x"c0",x"fe"),
  1526 => (x"87",x"c7",x"c9",x"49"),
  1527 => (x"c6",x"02",x"98",x"70"),
  1528 => (x"ea",x"fa",x"c1",x"87"),
  1529 => (x"c1",x"50",x"c1",x"48"),
  1530 => (x"bf",x"97",x"ea",x"fa"),
  1531 => (x"87",x"e3",x"c0",x"05"),
  1532 => (x"bf",x"f3",x"fa",x"c1"),
  1533 => (x"99",x"66",x"d0",x"49"),
  1534 => (x"87",x"d6",x"ff",x"05"),
  1535 => (x"bf",x"eb",x"fa",x"c1"),
  1536 => (x"99",x"66",x"d4",x"49"),
  1537 => (x"87",x"ca",x"ff",x"05"),
  1538 => (x"ed",x"e3",x"49",x"73"),
  1539 => (x"05",x"98",x"70",x"87"),
  1540 => (x"74",x"87",x"ff",x"fe"),
  1541 => (x"87",x"dc",x"fb",x"48"),
  1542 => (x"5c",x"5b",x"5e",x"0e"),
  1543 => (x"86",x"f4",x"0e",x"5d"),
  1544 => (x"ec",x"4c",x"4d",x"c0"),
  1545 => (x"a6",x"c4",x"7e",x"bf"),
  1546 => (x"f7",x"fa",x"c1",x"48"),
  1547 => (x"1e",x"c1",x"78",x"bf"),
  1548 => (x"49",x"c7",x"1e",x"c0"),
  1549 => (x"c8",x"87",x"cd",x"fd"),
  1550 => (x"02",x"98",x"70",x"86"),
  1551 => (x"49",x"ff",x"87",x"cd"),
  1552 => (x"c1",x"87",x"cc",x"fb"),
  1553 => (x"f1",x"e2",x"49",x"da"),
  1554 => (x"c1",x"4d",x"c1",x"87"),
  1555 => (x"bf",x"97",x"ea",x"fa"),
  1556 => (x"c7",x"87",x"c3",x"02"),
  1557 => (x"fa",x"c1",x"87",x"e6"),
  1558 => (x"c1",x"4b",x"bf",x"ef"),
  1559 => (x"05",x"bf",x"cf",x"e8"),
  1560 => (x"c3",x"87",x"e9",x"c0"),
  1561 => (x"d1",x"e2",x"49",x"fd"),
  1562 => (x"49",x"fa",x"c3",x"87"),
  1563 => (x"73",x"87",x"cb",x"e2"),
  1564 => (x"99",x"ff",x"c3",x"49"),
  1565 => (x"49",x"c0",x"1e",x"71"),
  1566 => (x"73",x"87",x"ce",x"fb"),
  1567 => (x"29",x"b7",x"c8",x"49"),
  1568 => (x"49",x"c1",x"1e",x"71"),
  1569 => (x"c8",x"87",x"c2",x"fb"),
  1570 => (x"87",x"fa",x"c5",x"86"),
  1571 => (x"bf",x"f3",x"fa",x"c1"),
  1572 => (x"dd",x"02",x"9b",x"4b"),
  1573 => (x"cb",x"e8",x"c1",x"87"),
  1574 => (x"c6",x"c6",x"49",x"bf"),
  1575 => (x"05",x"98",x"70",x"87"),
  1576 => (x"4b",x"c0",x"87",x"c4"),
  1577 => (x"e0",x"c2",x"87",x"d2"),
  1578 => (x"87",x"eb",x"c5",x"49"),
  1579 => (x"58",x"cf",x"e8",x"c1"),
  1580 => (x"e8",x"c1",x"87",x"c6"),
  1581 => (x"78",x"c0",x"48",x"cb"),
  1582 => (x"99",x"c2",x"49",x"73"),
  1583 => (x"c3",x"87",x"cd",x"05"),
  1584 => (x"f5",x"e0",x"49",x"eb"),
  1585 => (x"c2",x"49",x"70",x"87"),
  1586 => (x"87",x"c2",x"02",x"99"),
  1587 => (x"49",x"73",x"4c",x"fb"),
  1588 => (x"cd",x"05",x"99",x"c1"),
  1589 => (x"49",x"f4",x"c3",x"87"),
  1590 => (x"70",x"87",x"df",x"e0"),
  1591 => (x"02",x"99",x"c2",x"49"),
  1592 => (x"4c",x"fa",x"87",x"c2"),
  1593 => (x"99",x"c8",x"49",x"73"),
  1594 => (x"c3",x"87",x"cd",x"05"),
  1595 => (x"c9",x"e0",x"49",x"f5"),
  1596 => (x"c2",x"49",x"70",x"87"),
  1597 => (x"87",x"d4",x"02",x"99"),
  1598 => (x"bf",x"fb",x"fa",x"c1"),
  1599 => (x"48",x"87",x"c9",x"02"),
  1600 => (x"fa",x"c1",x"88",x"c1"),
  1601 => (x"87",x"c2",x"58",x"ff"),
  1602 => (x"4d",x"c1",x"4c",x"ff"),
  1603 => (x"99",x"c4",x"49",x"73"),
  1604 => (x"c3",x"87",x"ce",x"05"),
  1605 => (x"df",x"ff",x"49",x"f2"),
  1606 => (x"49",x"70",x"87",x"e0"),
  1607 => (x"db",x"02",x"99",x"c2"),
  1608 => (x"fb",x"fa",x"c1",x"87"),
  1609 => (x"c7",x"48",x"7e",x"bf"),
  1610 => (x"cb",x"03",x"a8",x"b7"),
  1611 => (x"c1",x"48",x"6e",x"87"),
  1612 => (x"ff",x"fa",x"c1",x"80"),
  1613 => (x"87",x"c2",x"c0",x"58"),
  1614 => (x"4d",x"c1",x"4c",x"fe"),
  1615 => (x"ff",x"49",x"fd",x"c3"),
  1616 => (x"70",x"87",x"f7",x"de"),
  1617 => (x"02",x"99",x"c2",x"49"),
  1618 => (x"fa",x"c1",x"87",x"d5"),
  1619 => (x"c0",x"02",x"bf",x"fb"),
  1620 => (x"fa",x"c1",x"87",x"c9"),
  1621 => (x"78",x"c0",x"48",x"fb"),
  1622 => (x"fd",x"87",x"c2",x"c0"),
  1623 => (x"c3",x"4d",x"c1",x"4c"),
  1624 => (x"de",x"ff",x"49",x"fa"),
  1625 => (x"49",x"70",x"87",x"d4"),
  1626 => (x"d9",x"02",x"99",x"c2"),
  1627 => (x"fb",x"fa",x"c1",x"87"),
  1628 => (x"b7",x"c7",x"48",x"bf"),
  1629 => (x"c9",x"c0",x"03",x"a8"),
  1630 => (x"fb",x"fa",x"c1",x"87"),
  1631 => (x"c0",x"78",x"c7",x"48"),
  1632 => (x"4c",x"fc",x"87",x"c2"),
  1633 => (x"b7",x"c0",x"4d",x"c1"),
  1634 => (x"d1",x"c0",x"03",x"ac"),
  1635 => (x"4a",x"66",x"c4",x"87"),
  1636 => (x"6a",x"82",x"d8",x"c1"),
  1637 => (x"87",x"c6",x"c0",x"02"),
  1638 => (x"49",x"74",x"4b",x"6a"),
  1639 => (x"1e",x"c0",x"0f",x"73"),
  1640 => (x"c1",x"1e",x"f0",x"c3"),
  1641 => (x"db",x"f7",x"49",x"da"),
  1642 => (x"70",x"86",x"c8",x"87"),
  1643 => (x"e2",x"c0",x"02",x"98"),
  1644 => (x"48",x"a6",x"c8",x"87"),
  1645 => (x"bf",x"fb",x"fa",x"c1"),
  1646 => (x"49",x"66",x"c8",x"78"),
  1647 => (x"66",x"c4",x"91",x"cb"),
  1648 => (x"70",x"80",x"71",x"48"),
  1649 => (x"02",x"bf",x"6e",x"7e"),
  1650 => (x"6e",x"87",x"c8",x"c0"),
  1651 => (x"66",x"c8",x"4b",x"bf"),
  1652 => (x"75",x"0f",x"73",x"49"),
  1653 => (x"c8",x"c0",x"02",x"9d"),
  1654 => (x"fb",x"fa",x"c1",x"87"),
  1655 => (x"c9",x"f3",x"49",x"bf"),
  1656 => (x"d3",x"e8",x"c1",x"87"),
  1657 => (x"dd",x"c0",x"02",x"bf"),
  1658 => (x"f6",x"c0",x"49",x"87"),
  1659 => (x"02",x"98",x"70",x"87"),
  1660 => (x"c1",x"87",x"d3",x"c0"),
  1661 => (x"49",x"bf",x"fb",x"fa"),
  1662 => (x"c0",x"87",x"ef",x"f2"),
  1663 => (x"87",x"cf",x"f4",x"49"),
  1664 => (x"48",x"d3",x"e8",x"c1"),
  1665 => (x"8e",x"f4",x"78",x"c0"),
  1666 => (x"00",x"87",x"e9",x"f3"),
  1667 => (x"00",x"00",x"00",x"00"),
  1668 => (x"00",x"00",x"00",x"00"),
  1669 => (x"1e",x"00",x"00",x"00"),
  1670 => (x"c8",x"ff",x"4a",x"71"),
  1671 => (x"a1",x"72",x"49",x"bf"),
  1672 => (x"1e",x"4f",x"26",x"48"),
  1673 => (x"89",x"bf",x"c8",x"ff"),
  1674 => (x"c0",x"c0",x"c0",x"c2"),
  1675 => (x"01",x"a9",x"c0",x"c0"),
  1676 => (x"4a",x"c0",x"87",x"c4"),
  1677 => (x"4a",x"c1",x"87",x"c2"),
  1678 => (x"4f",x"26",x"48",x"72"),
  1679 => (x"e5",x"e9",x"c1",x"1e"),
  1680 => (x"b9",x"c1",x"49",x"bf"),
  1681 => (x"59",x"e9",x"e9",x"c1"),
  1682 => (x"c3",x"48",x"d4",x"ff"),
  1683 => (x"d0",x"ff",x"78",x"ff"),
  1684 => (x"78",x"e1",x"c0",x"48"),
  1685 => (x"c1",x"48",x"d4",x"ff"),
  1686 => (x"71",x"31",x"c4",x"78"),
  1687 => (x"48",x"d0",x"ff",x"78"),
  1688 => (x"26",x"78",x"e0",x"c0"),
  1689 => (x"00",x"00",x"00",x"4f"),
  1690 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

