//-------------------------------------------------------------------------------------------------
module spi
//-------------------------------------------------------------------------------------------------
(
	input  wire      clock,
	input  wire      ce,
	input  wire      io,
	input  wire[7:0] d,
	output reg [7:0] q,
	output wire      ck,
	output wire      mosi,
	input  wire      miso
);
//-------------------------------------------------------------------------------------------------

reg[7:0] sd;
reg[4:0] count = 5'b10000;

always @(posedge clock) if(ce)
	if(count[4]) begin
		if(io) begin
			q <= sd;
			sd <= d;
			count <= 5'd0;
		end
	end
	else begin
		count <= count+5'd1;
		if(count[0]) sd <= { sd[6:0], miso };
	end

//-------------------------------------------------------------------------------------------------

assign ck = count[0];
assign mosi = sd[7];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
