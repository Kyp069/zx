//-------------------------------------------------------------------------------------------------
// x-axis  64479 FBDF xxxxx011 xx0xxxxx
// y-axis  65503 FFDF xxxxx111 xx0xxxxx
// 
// buttons 64223 FADF xxxxxx10 xx0xxxxx
// 
// D[0] = right button
// D[1] = left button
// D[2] = middle button
// D[3] = floating bus
// D[7:4] = wheel counter
//-------------------------------------------------------------------------------------------------
module mouse
//-------------------------------------------------------------------------------------------------
(
);
//-------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
